* NGSPICE file created from controller_core.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyd_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyd_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyd_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyd_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_2 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

.subckt controller_core clock clock_out[0] clock_out[1] clock_out[2] clock_out[3]
+ clock_out[4] clock_out[5] clock_out[6] clock_out[7] clock_out[8] clock_out[9] col_select_left[0]
+ col_select_left[1] col_select_left[2] col_select_left[3] col_select_left[4] col_select_left[5]
+ col_select_right[0] col_select_right[1] col_select_right[2] col_select_right[3]
+ col_select_right[4] col_select_right[5] data_out_left[0] data_out_left[10] data_out_left[11]
+ data_out_left[12] data_out_left[13] data_out_left[14] data_out_left[15] data_out_left[1]
+ data_out_left[2] data_out_left[3] data_out_left[4] data_out_left[5] data_out_left[6]
+ data_out_left[7] data_out_left[8] data_out_left[9] data_out_right[0] data_out_right[10]
+ data_out_right[11] data_out_right[12] data_out_right[13] data_out_right[14] data_out_right[15]
+ data_out_right[1] data_out_right[2] data_out_right[3] data_out_right[4] data_out_right[5]
+ data_out_right[6] data_out_right[7] data_out_right[8] data_out_right[9] inverter_select[0]
+ inverter_select[1] inverter_select[2] inverter_select[3] inverter_select[4] inverter_select[5]
+ inverter_select[6] inverter_select[7] inverter_select[8] inverter_select[9] io_control_trigger_in
+ io_control_trigger_oeb io_driver_io_oeb[0] io_driver_io_oeb[10] io_driver_io_oeb[11]
+ io_driver_io_oeb[12] io_driver_io_oeb[13] io_driver_io_oeb[14] io_driver_io_oeb[15]
+ io_driver_io_oeb[16] io_driver_io_oeb[17] io_driver_io_oeb[18] io_driver_io_oeb[19]
+ io_driver_io_oeb[1] io_driver_io_oeb[2] io_driver_io_oeb[3] io_driver_io_oeb[4]
+ io_driver_io_oeb[5] io_driver_io_oeb[6] io_driver_io_oeb[7] io_driver_io_oeb[8]
+ io_driver_io_oeb[9] io_latch_data_in io_latch_data_oeb io_reset_n_in io_reset_n_oeb
+ io_update_cycle_complete_oeb io_update_cycle_complete_out la_data_in[0] la_data_in[10]
+ la_data_in[11] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16]
+ la_data_in[17] la_data_in[1] la_data_in[2] la_data_in[3] la_data_in[4] la_data_in[5]
+ la_data_in[6] la_data_in[7] la_data_in[8] la_data_in[9] la_oenb[0] la_oenb[10] la_oenb[11]
+ la_oenb[12] la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[1]
+ la_oenb[2] la_oenb[3] la_oenb[4] la_oenb[5] la_oenb[6] la_oenb[7] la_oenb[8] la_oenb[9]
+ mem_address_left[0] mem_address_left[1] mem_address_left[2] mem_address_left[3]
+ mem_address_left[4] mem_address_left[5] mem_address_left[6] mem_address_left[7]
+ mem_address_left[8] mem_address_left[9] mem_address_right[0] mem_address_right[1]
+ mem_address_right[2] mem_address_right[3] mem_address_right[4] mem_address_right[5]
+ mem_address_right[6] mem_address_right[7] mem_address_right[8] mem_address_right[9]
+ mem_write_n[0] mem_write_n[1] mem_write_n[2] mem_write_n[3] mem_write_n[4] mem_write_n[5]
+ mem_write_n[6] mem_write_n[7] mem_write_n[8] mem_write_n[9] output_active_left output_active_right
+ row_col_select[0] row_col_select[1] row_col_select[2] row_col_select[3] row_col_select[4]
+ row_col_select[5] row_col_select[6] row_col_select[7] row_col_select[8] row_col_select[9]
+ row_select_left[0] row_select_left[1] row_select_left[2] row_select_left[3] row_select_left[4]
+ row_select_left[5] row_select_right[0] row_select_right[1] row_select_right[2] row_select_right[3]
+ row_select_right[4] row_select_right[5] spi_data[0] spi_data[10] spi_data[11] spi_data[12]
+ spi_data[13] spi_data[14] spi_data[15] spi_data[16] spi_data[17] spi_data[18] spi_data[19]
+ spi_data[1] spi_data[20] spi_data[21] spi_data[22] spi_data[23] spi_data[24] spi_data[25]
+ spi_data[26] spi_data[27] spi_data[28] spi_data[29] spi_data[2] spi_data[30] spi_data[31]
+ spi_data[3] spi_data[4] spi_data[5] spi_data[6] spi_data[7] spi_data[8] spi_data[9]
+ spi_data_clock vdd vss
XFILLER_45_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3155_ spi_data_crossing\[18\].A clknet_leaf_5_clock spi_data_crossing\[18\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3086_ _0220_ clknet_leaf_29_clock u1.timer\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2106_ _0404_ _0495_ _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2037_ _0448_ _0076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2246__A3 _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2939_ _0081_ clknet_leaf_4_clock u1.ordering_complete\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1757__A2 _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2706__A1 _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3171__D spi_data_crossing\[26\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1479__I u1.ordering_complete\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1445__A1 _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2642__B1 _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1996__A2 _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2796__I1 _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2712__A4 _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2476__A3 _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3005__CLK clknet_leaf_12_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2724_ _0968_ _0973_ _0974_ _0237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2655_ u1.ccr1\[18\] _0920_ _0921_ _0922_ _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__3155__CLK clknet_leaf_5_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1606_ _1223_ _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2164__A2 _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2586_ u0.cmd\[29\] _0864_ _0865_ spi_data_crossing\[29\].data_sync _0867_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1537_ _1157_ u0.latch_cmd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1468_ _1072_ _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3207_ _0277_ clknet_leaf_35_clock net159 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3138_ net41 net230 spi_data_crossing\[10\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2683__I _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3069_ _0210_ clknet_leaf_9_clock u1.row_sel\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2794__S _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2458__A3 _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1418__A1 _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2091__A1 net220 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3028__CLK clknet_leaf_24_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1969__A2 _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1937__I net223 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2440_ _0759_ _0168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_45_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2371_ _1100_ _0694_ _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1672__I u1.timer\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2621__A3 _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2707_ _1311_ _0961_ _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_12_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2137__A2 _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2638_ u1.ccr1\[11\] _1269_ u1.ccr1\[10\] _1268_ _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_12_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2569_ _0856_ _0200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1582__I u1.ccr1\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input36_I la_oenb[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1648__A1 _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3302__I net168 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1820__A1 _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_15_clock_I clknet_2_3__leaf_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2300__A2 _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2029__S _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1940_ _0353_ _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1871_ net226 _0332_ _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_fanout223_I u0.cmd\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2119__A2 _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2423_ _0744_ _0166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1878__A1 u1.col_sel\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2354_ _1103_ _0683_ _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2285_ u1.ordering_timer\[3\] _0602_ _0605_ _0623_ _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_38_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2358__A2 _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1869__A1 u0.timer_enable vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2201__I _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2294__A1 _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2597__A2 _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1487__I u1.ordering_complete\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2860__CLK clknet_leaf_9_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3216__CLK clknet_leaf_17_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2070_ _0455_ _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_35_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2972_ _0114_ clknet_leaf_9_clock u1.row_limit\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1923_ _1329_ _0360_ _0372_ _0038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1854_ u1.col_sel\[1\] _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_19_clock clknet_2_3__leaf_clock clknet_leaf_19_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1785_ _1212_ _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2060__I1 u1.ordering_complete\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2406_ u1.ordering_complete\[18\] _0714_ _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2337_ _0669_ _0155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2268_ _0608_ _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_38_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2276__A1 _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2199_ _0551_ _0135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2883__CLK clknet_leaf_9_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3239__CLK clknet_leaf_7_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2200__A1 u0.cmd\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3174__D net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold41 u1.row_col_select\[2\] net283 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold30 latch_data_sync\[0\] net272 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold52 u1.col_sel\[4\] net294 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_25_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1490__A2 _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1778__B1 _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2042__S _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2042__I1 _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1570_ u1.timer\[6\] _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3240_ net258 clknet_leaf_7_clock net168 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3171_ spi_data_crossing\[26\].A clknet_leaf_7_clock spi_data_crossing\[26\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2122_ _0478_ u1.ordering_complete\[25\] _0489_ _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_48_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2053_ _0356_ _0458_ _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_19_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2217__S _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1481__A2 u1.ordering_complete\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2955_ _0097_ clknet_leaf_3_clock u1.ordering_complete\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2886_ _0020_ clknet_leaf_8_clock u0.mem_write_n\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1906_ _0359_ _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1837_ _0302_ _0303_ _0305_ _0018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_15_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1768_ _1256_ u1.ccr0\[15\] _1306_ _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_46_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1699_ _1302_ _1308_ _1309_ _1315_ _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XTAP_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2497__A1 _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1590__I u1.timer\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3310__I net207 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output105_I net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3061__CLK clknet_leaf_7_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3169__D spi_data_crossing\[25\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2421__A1 _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput75 net75 clock_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
XFILLER_1_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput86 net86 col_select_left[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_49_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput97 net97 data_out_left[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__2488__A1 _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2660__A1 u1.ccr1\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2412__A1 u1.ordering_timer\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2740_ _0983_ _0984_ _0985_ _0242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2671_ _0933_ _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1622_ u1.ccr1\[18\] u1.timer\[18\] _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1553_ u1.timer\[31\] _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1484_ u1.ordering_timer\[9\] _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_28_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3223_ net265 clknet_leaf_17_clock net136 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3154_ net49 net235 spi_data_crossing\[18\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2105_ _0491_ _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3085_ _0219_ clknet_leaf_35_clock net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2036_ u1.ccr1\[28\] _0447_ _0443_ _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3084__CLK clknet_leaf_4_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2651__A1 _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2938_ _0080_ clknet_leaf_12_clock u1.ordering_complete\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2869_ _0026_ clknet_leaf_10_clock u1.col_sel\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2921__CLK clknet_leaf_29_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input66_I spi_data[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2706__A2 _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1534__B _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2190__I0 _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_2_1__f_clock_I clknet_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2181__I0 _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2944__CLK clknet_leaf_19_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2723_ _0282_ u1.timer\[16\] _0970_ _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__1739__A3 _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2654_ _0434_ u1.timer\[19\] _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2585_ _0866_ _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1605_ u1.timer\[20\] _1223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1536_ _1156_ u0.u11.impulse_gen\[1\] _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_47_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1467_ _1088_ u1.ordering_complete\[25\] _1091_ _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_41_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3206_ _0276_ clknet_leaf_29_clock u1.ccr0\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3137_ spi_data_crossing\[9\].A clknet_leaf_0_clock spi_data_crossing\[9\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3068_ _0023_ clknet_leaf_4_clock u1.output_active vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2624__A1 _0890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2019_ _0438_ _0068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3182__D _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2615__A1 u1.row_sel\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1418__A2 u0.cmd\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2967__CLK clknet_leaf_23_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_11_clock_I clknet_2_1__leaf_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1953__I u0.cmd\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2370_ u1.ordering_timer\[14\] _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1657__A2 _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3122__CLK net229 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2706_ _0958_ _0961_ _0962_ _0231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
Xoutput210 net210 row_select_right[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_2637_ _0905_ net38 _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_12_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2568_ u0.cmd\[22\] _0852_ _0853_ spi_data_crossing\[22\].data_sync _0856_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1519_ _1070_ _1095_ _1120_ _1143_ _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__1896__A2 _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2499_ u1.ordering_timer\[31\] _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2145__I0 _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input29_I la_oenb[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3177__D spi_data_crossing\[29\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1959__I0 u1.ccr1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output97_I net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3145__CLK clknet_leaf_1_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1870_ net226 _0332_ _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_30_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1683__I u1.timer\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2422_ u1.ordering_timer\[20\] _0719_ _0733_ _0743_ _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2353_ _0675_ _0677_ _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2284_ _0613_ _0621_ _0622_ _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1802__A2 _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1999_ _0388_ _0398_ _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1566__A1 u1.ccr1\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3018__CLK clknet_leaf_13_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1869__A2 _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2818__A1 u0.cmd\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2046__A2 u0.cmd\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1557__A1 _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2285__A2 _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2971_ _0113_ clknet_leaf_11_clock u1.row_limit\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1922_ _0370_ _0371_ _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1853_ u1.col_sel\[2\] _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1784_ _1292_ _1374_ _1400_ _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2405_ _0728_ _0723_ _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2336_ u1.ordering_timer\[9\] _0655_ _0662_ _0668_ _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1720__A1 _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2267_ _0607_ _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2198_ _0478_ u1.inverter_select\[9\] _0539_ _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_1_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3308__I net205 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold31 u1.row_col_select\[1\] net273 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold20 u1.inverter_select\[4\] net262 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_0_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold42 u1.row_col_select\[7\] net284 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold53 u1.col_sel\[1\] net295 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XANTENNA__3190__D _0260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1950__A1 _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1961__I u0.cmd\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3170_ net58 net237 spi_data_crossing\[26\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2121_ _0504_ _0104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2052_ _1133_ _0457_ _0459_ _0080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_48_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2502__I0 u1.ordering_complete\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2954_ _0096_ clknet_leaf_3_clock u1.ordering_complete\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2885_ _0019_ clknet_leaf_8_clock u0.mem_write_n\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1905_ _0352_ _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1836_ _0301_ _0305_ _0017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1767_ _1302_ _1308_ _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_1_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1941__A1 net222 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1698_ _1312_ _1314_ _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2497__A2 _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2319_ _0653_ _0153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3299_ net165 net175 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2850__CLK clknet_leaf_15_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input11_I la_data_in[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3206__CLK clknet_leaf_29_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2143__S _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3185__D _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput76 net76 clock_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
XFILLER_27_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput98 net98 data_out_left[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput87 net87 col_select_left[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_27_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2488__A2 _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_18_clock clknet_2_3__leaf_clock clknet_leaf_18_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_29_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1999__A1 _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2117__I _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2412__A2 _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2670_ _0935_ _0936_ _0221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1620__B1 u1.ccr1\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1621_ u1.ccr1\[19\] u1.timer\[19\] _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1552_ u1.ccr1\[25\] _1164_ u1.ccr1\[24\] _1166_ _1169_ _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XANTENNA__1923__A1 _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1483_ _1099_ _1102_ _1107_ _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2787__I _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3222_ net278 clknet_leaf_18_clock net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2873__CLK clknet_leaf_16_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3153_ spi_data_crossing\[17\].A clknet_leaf_5_clock spi_data_crossing\[17\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2479__A2 _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input3_I io_reset_n_in vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2104_ _1061_ _0490_ _0494_ _0097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3084_ _0010_ clknet_leaf_4_clock u0.run_state\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2736__B _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3229__CLK clknet_leaf_18_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2035_ net222 _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1866__I _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2937_ _0079_ clknet_leaf_0_clock u1.ccr1\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2868_ _0025_ clknet_leaf_11_clock u1.col_sel\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2167__A1 _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1819_ u0.cmd\[30\] _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2799_ _0409_ _1021_ _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_2_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input59_I spi_data[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2896__CLK clknet_leaf_2_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2330__A1 _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2181__I1 u1.inverter_select\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2633__A2 latch_data vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1686__I u1.timer\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2397__A1 _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2722_ _0283_ _0971_ _0282_ _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_34_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2653_ _1241_ _1238_ _1242_ _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2584_ u0.cmd\[28\] _0864_ _0865_ spi_data_crossing\[28\].data_sync _0866_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_12_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1604_ _1202_ _1211_ _1221_ _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1535_ u0.u11.impulse_gen\[0\] _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1466_ u1.ordering_timer\[24\] _1086_ _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3205_ _0275_ clknet_leaf_23_clock u1.ccr0\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3051__CLK clknet_leaf_1_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3136_ net71 net230 spi_data_crossing\[9\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3067_ _0209_ clknet_leaf_6_clock u0.cmd\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2018_ u1.ccr1\[20\] _0366_ _0432_ _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_35_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output165_I net165 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2560__B2 spi_data_crossing\[19\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2560__A1 net218 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2615__A2 _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1418__A3 _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3074__CLK clknet_leaf_10_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2303__A1 u1.ordering_complete\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2911__CLK clknet_leaf_24_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2705_ _1272_ _0959_ _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xoutput200 net200 row_col_select[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_2636_ net20 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1593__A2 _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput211 net211 row_select_right[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_2567_ _0855_ _0199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2542__A1 _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1518_ _1132_ _1135_ _1137_ _1142_ _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_2498_ _0565_ _0602_ _0808_ _0809_ _0176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1449_ u1.ordering_timer\[31\] _1073_ _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2145__I1 u1.row_limit\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3119_ spi_data_crossing\[0\].A clknet_leaf_35_clock spi_data_crossing\[0\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3097__CLK clknet_leaf_26_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1959__I1 _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1990__S _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2934__CLK clknet_leaf_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1964__I _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2772__A1 _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2421_ _0734_ _0741_ _0742_ _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2524__A1 _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2352_ _0626_ _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2524__B2 spi_data_crossing\[5\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2283_ u1.ordering_complete\[3\] _0597_ _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2035__I net222 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2063__I0 _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1998_ _1263_ _0421_ _0424_ _0061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2763__A1 _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1566__A2 _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2619_ u1.row_sel\[2\] u1.row_sel\[1\] _0892_ _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__2957__CLK clknet_leaf_3_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input41_I spi_data[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2046__A3 u0.cmd\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3188__D _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3112__CLK clknet_leaf_34_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2970_ _0112_ clknet_leaf_12_clock u1.row_limit\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1921_ _0353_ _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1852_ _0313_ u1.col_limit\[3\] _0314_ u1.col_limit\[4\] _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__2745__A1 _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1783_ _1362_ _1393_ _1399_ _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2404_ _1065_ _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_44_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2335_ _0643_ _0666_ _0667_ _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_38_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2266_ _0595_ _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2197_ _0550_ _0134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2036__I0 u1.ccr1\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2736__A1 _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3135__CLK clknet_leaf_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold32 u1.row_col_select\[3\] net274 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold10 u0.mem_write_n\[0\] net252 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold21 u1.row_col_select\[4\] net263 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold43 u0.cmd\[24\] net285 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_28_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1778__A2 _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2727__A1 _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2403__I _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2120_ _0476_ u1.ordering_complete\[24\] _0498_ _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2051_ _0345_ _0458_ _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_19_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2663__B1 _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2953_ _0095_ clknet_leaf_3_clock u1.ordering_complete\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3008__CLK clknet_leaf_14_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1904_ _0358_ _0033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2884_ _0018_ clknet_leaf_8_clock u0.mem_write_n\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1835_ _0298_ _0305_ _0016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1766_ _1313_ _1382_ _1312_ _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_15_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1697_ _1267_ u1.ccr0\[8\] _1313_ _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2318_ _0648_ _0627_ _0635_ _0652_ _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3298_ net164 net174 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2249_ _1080_ _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2223__I _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2709__A1 _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput88 net88 col_select_left[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput77 net77 clock_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
Xoutput99 net99 data_out_left[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_27_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2488__A3 _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1620__B2 _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1620__A1 u1.ccr1\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1620_ u1.ccr1\[17\] _1236_ u1.ccr1\[16\] _1237_ _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__2176__A2 _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1551_ u1.ccr1\[30\] _1167_ u1.ccr1\[29\] _1168_ _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__1923__A2 _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1482_ _1103_ u1.ordering_complete\[12\] _1105_ _1106_ _1107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3221_ net282 clknet_leaf_17_clock net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3152_ net48 net234 spi_data_crossing\[17\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2103_ _0356_ _0492_ _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3083_ _0009_ clknet_leaf_4_clock u0.run_state\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2736__C _0982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2034_ _1176_ _0436_ _0446_ _0075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2936_ _0078_ clknet_leaf_0_clock u1.ccr1\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2867_ _0024_ clknet_leaf_32_clock net160 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1818_ _0294_ _0005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2167__A2 _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2798_ _1012_ _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1749_ _1363_ u1.ccr0\[1\] _1365_ _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output110_I net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1602__A1 _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2094__A1 _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2128__I _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1841__A1 _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1967__I _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout239_I net240 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2397__A2 _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2721_ _1279_ _0932_ _0971_ _0283_ _0972_ _0236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_12_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2652_ _0434_ _1318_ _1321_ _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2840__CLK clknet_leaf_15_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2583_ _0846_ _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1603_ _1212_ _1216_ _1217_ _1220_ _1221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__2798__I _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1534_ _1153_ _1154_ _1155_ _0006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2990__CLK clknet_leaf_17_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1465_ _1085_ _1086_ _1089_ _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3204_ _0274_ clknet_leaf_23_clock u1.ccr0\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3135_ spi_data_crossing\[8\].A clknet_leaf_0_clock spi_data_crossing\[8\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3066_ _0208_ clknet_leaf_6_clock u0.cmd\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2085__A1 net223 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2017_ _0434_ _0435_ _0437_ _0067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_24_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2919_ _0061_ clknet_leaf_27_clock u1.ccr1\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_17_clock clknet_2_3__leaf_clock clknet_leaf_17_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_input71_I spi_data[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1787__I _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2863__CLK clknet_leaf_4_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3219__CLK clknet_leaf_17_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2000__A1 _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2303__A2 _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2704_ _1272_ u1.timer\[10\] _0950_ _0955_ _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
Xoutput201 net201 row_col_select[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_2635_ _1156_ _0815_ _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_12_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2790__A2 _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput212 net212 row_select_right[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_47_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2566_ u0.cmd\[21\] _0852_ _0853_ spi_data_crossing\[21\].data_sync _0855_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1517_ _1139_ u1.ordering_complete\[0\] _1140_ _1141_ _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_2497_ _1082_ _0716_ _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1448_ u1.ordering_complete\[31\] _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3118_ net40 net227 spi_data_crossing\[0\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3049_ _0191_ clknet_leaf_4_clock u0.cmd\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2886__CLK clknet_leaf_8_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1805__A1 _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3041__CLK clknet_leaf_4_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2420_ u1.ordering_complete\[20\] _0687_ _0742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3191__CLK clknet_leaf_23_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2351_ _0681_ _0157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1980__I _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2282_ u1.ordering_timer\[3\] _0614_ _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_9_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2460__A1 _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1997_ net221 _0418_ _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2063__I1 u1.ordering_complete\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2618_ _0891_ _0894_ _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1890__I _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2549_ _0843_ _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_47_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input34_I la_oenb[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2279__A1 _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2000__B _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3064__CLK clknet_leaf_6_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2754__A2 _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2901__CLK clknet_leaf_34_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1493__A2 _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1920_ u0.cmd\[6\] _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1851_ u1.col_sel\[4\] _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_42_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout221_I u0.cmd\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1782_ _1171_ u1.ccr0\[31\] _1354_ _1398_ _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_7_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2403_ _0727_ _0163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_48_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2334_ _1110_ _0658_ _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2265_ _1138_ _0599_ _0606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2196_ _0476_ u1.inverter_select\[8\] _0539_ _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_38_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3087__CLK clknet_leaf_29_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2808__I0 u1.ccr0\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1641__C1 u1.ccr1\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2924__CLK clknet_leaf_3_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2036__I1 _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold22 u1.row_col_select\[6\] net264 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold11 u1.inverter_select\[3\] net253 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold33 u1.inverter_select\[2\] net275 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold44 u0.cmd\[25\] net286 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_25_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold42_I u1.row_col_select\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2360__B1 _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2050_ _0456_ _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2663__A1 _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2947__CLK clknet_leaf_20_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2415__A1 u1.ordering_complete\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2952_ _0094_ clknet_leaf_3_clock u1.ordering_complete\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1903_ u1.ccr0\[17\] _0357_ _0354_ _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2883_ _0017_ clknet_leaf_9_clock u0.mem_write_n\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1834_ _0304_ u0.cmd\[29\] _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_11_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2018__I1 _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1765_ _1294_ _1297_ _1299_ _1309_ _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_11_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1696_ _1262_ _1310_ _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3297_ net163 net173 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2317_ _0643_ _0650_ _0651_ _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2248_ _1084_ _0589_ _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_39_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2485__B _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2179_ _0346_ u1.inverter_select\[0\] _0540_ _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_38_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2406__A1 u1.ordering_complete\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3102__CLK clknet_leaf_28_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2709__A2 _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1564__B _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3252__CLK clknet_leaf_9_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput89 net89 col_select_right[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput78 net78 clock_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
XFILLER_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2342__B1 _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2488__A4 _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1696__A2 _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1620__A2 _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1550_ u1.timer\[29\] _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1481_ _1101_ u1.ordering_complete\[13\] _1103_ u1.ordering_complete\[12\] _1106_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3220_ net281 clknet_leaf_17_clock net133 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3151_ spi_data_crossing\[16\].A clknet_leaf_5_clock spi_data_crossing\[16\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2102_ _1060_ _0490_ _0493_ _0096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1931__I0 u1.ccr0\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3082_ _0008_ clknet_leaf_4_clock u0.run_state\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2033_ _0382_ _0428_ _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3125__CLK clknet_leaf_36_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2935_ _0077_ clknet_leaf_0_clock u1.ccr1\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2324__I _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2866_ net259 clknet_leaf_34_clock reset_n_sync\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1817_ _1153_ u0.run_state\[0\] _1155_ _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_11_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2797_ _1020_ _0264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1748_ _1363_ u1.ccr0\[1\] u1.ccr0\[0\] _1364_ _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1679_ u1.ccr0\[10\] _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2627__A1 _0890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output103_I net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2618__A1 _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2094__A2 _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2633__A4 _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2720_ _0283_ _0971_ _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2651_ _1227_ _1231_ _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2080__S _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1602_ _1218_ _1219_ _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2582_ _0844_ _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1533_ _1040_ u0.cmd\[30\] _1042_ _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_1464_ _1087_ u1.ordering_complete\[26\] _1088_ u1.ordering_complete\[25\] _1089_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3203_ _0273_ clknet_leaf_23_clock u1.ccr0\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_0_clock clock clknet_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3134_ net70 net230 spi_data_crossing\[8\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2609__B2 net216 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3065_ _0207_ clknet_leaf_6_clock u0.cmd\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2016_ _0407_ _0436_ _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1832__A2 _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2918_ _0060_ clknet_leaf_27_clock u1.ccr1\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2849_ net289 clknet_leaf_16_clock net106 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1893__I net218 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input64_I spi_data[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2229__I _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2673__B _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1823__A2 u0.cmd\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2000__A2 _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2703_ _0958_ _0959_ _0960_ _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_12_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2634_ _0904_ _0217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput213 net213 row_select_right[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput202 net202 row_col_select[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_2565_ _0854_ _0198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1516_ _1136_ u1.ordering_complete\[2\] _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2496_ _0804_ _0807_ _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_4_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1447_ u1.ordering_timer\[27\] _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2049__I _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3117_ _0251_ clknet_leaf_36_clock u1.timer\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3048_ _0190_ clknet_leaf_5_clock u0.cmd\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1805__A2 _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_2_0__f_clock_I clknet_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output170_I net170 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2834__D u1.row_sel\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2980__CLK clknet_leaf_14_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2350_ _0675_ _0655_ _0662_ _0680_ _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2281_ _0620_ _0148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_16_clock clknet_2_3__leaf_clock clknet_leaf_16_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_25_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2460__A2 _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1996_ _1261_ _0421_ _0423_ _0060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1971__A1 _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2617_ _0878_ _0892_ _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2548_ _0390_ _0838_ _0839_ spi_data_crossing\[15\].data_sync _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_47_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2479_ _0508_ _0711_ _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2853__CLK clknet_leaf_16_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input27_I la_oenb[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2507__I _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3209__CLK clknet_leaf_28_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2451__A2 _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output95_I net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1850_ u1.col_sel\[3\] _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_30_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1781_ _1360_ _1397_ _1398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2745__A3 _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2402_ _1068_ _0719_ _0691_ _0726_ _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2876__CLK clknet_leaf_6_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2333_ _0664_ _0665_ _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2264_ _0604_ _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2195_ _0549_ _0133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1469__B1 _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2681__A2 _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2808__I1 _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2062__I _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1979_ _1196_ _0403_ _0413_ _0053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1944__A1 _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold23 u1.inverter_select\[9\] net265 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold12 u0.cmd\[23\] net254 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold45 u1.row_col_select\[0\] net287 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold34 u1.row_sel\[5\] net276 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_28_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3031__CLK clknet_leaf_24_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3181__CLK clknet_leaf_7_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2424__A2 _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2173__S _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2899__CLK clknet_leaf_36_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1935__A1 _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2700__I _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_hold35_I u1.inverter_select\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2663__A2 _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2415__A2 _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2951_ _0093_ clknet_leaf_4_clock u1.ordering_complete\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1902_ _0356_ _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2882_ _0016_ clknet_leaf_8_clock u0.mem_write_n\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1833_ u0.cmd\[28\] _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_30_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1926__A1 _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1764_ _1377_ _1378_ _1380_ _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_7_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1695_ _1300_ _1301_ _1310_ _1311_ _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_48_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3054__CLK clknet_leaf_5_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3296_ net162 net172 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2316_ u1.ordering_complete\[7\] _0630_ _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2247_ u1.ordering_timer\[27\] _0508_ u1.ordering_timer\[26\] _0506_ _1089_ _1092_
+ _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_38_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2103__A1 _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2178_ _0539_ _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_25_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2406__A2 _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2590__A1 _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1564__C _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2520__I _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput79 net79 clock_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
XANTENNA__2342__A1 u1.ordering_timer\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3077__CLK clknet_leaf_4_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1480_ u1.ordering_timer\[15\] _1097_ u1.ordering_timer\[11\] _1104_ _1105_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3150_ net47 net234 spi_data_crossing\[16\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3081_ _0007_ clknet_leaf_4_clock u0.run_state\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2101_ _0345_ _0492_ _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1931__I1 _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3261__I clknet_leaf_10_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2914__CLK clknet_leaf_25_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2032_ _1178_ _0435_ _0445_ _0074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2934_ _0076_ clknet_leaf_0_clock u1.ccr1\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2865_ net270 clknet_leaf_33_clock reset_n_sync\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1816_ net37 _1144_ _0293_ _0001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_15_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2796_ u1.ccr0\[3\] _0364_ _1013_ _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1747_ _1207_ _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1678_ u1.timer\[10\] _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3279_ net110 net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2515__I _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2315__A1 _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2937__CLK clknet_leaf_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1841__A3 _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2650_ _1266_ _0908_ _0910_ _0917_ _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_8_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1601_ _1213_ u1.timer\[3\] _1219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3256__I clknet_leaf_9_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2581_ _0863_ _0205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2160__I _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2554__A1 _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1532_ u0.run_state\[0\] _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1463_ u1.ordering_timer\[25\] _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3202_ _0272_ clknet_leaf_23_clock u1.ccr0\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input1_I io_control_trigger_in vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3133_ spi_data_crossing\[7\].A clknet_leaf_5_clock spi_data_crossing\[7\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3064_ _0206_ clknet_leaf_6_clock u0.cmd\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2015_ _0427_ _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3242__CLK clknet_leaf_7_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2917_ _0059_ clknet_leaf_26_clock u1.ccr1\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2848_ net290 clknet_leaf_16_clock net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2070__I _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2779_ net5 _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input57_I spi_data[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_9_clock_I clknet_2_1__leaf_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2181__S _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2784__A1 _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1587__A2 _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2536__A1 _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2536__B2 spi_data_crossing\[10\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3115__CLK clknet_leaf_36_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2702_ _1295_ _0956_ _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_13_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2633_ latch_data_sync\[0\] latch_data latch_data_sync\[1\] _1042_ _0904_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__and4_1
Xoutput214 net214 row_select_right[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput203 net203 row_col_select[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_2564_ u0.cmd\[20\] _0852_ _0853_ spi_data_crossing\[20\].data_sync _0854_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1515_ u1.ordering_timer\[1\] _1134_ _1140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2495_ _1082_ _0801_ _0805_ _0806_ _0780_ _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_1446_ u1.ordering_timer\[28\] _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3116_ _0250_ clknet_leaf_36_clock u1.timer\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3047_ _0189_ clknet_leaf_1_clock u0.cmd\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1805__A3 u1.timer\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2065__I _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2066__I0 _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1569__A2 _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1813__I0 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2518__A1 _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2518__B2 spi_data_crossing\[3\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output163_I net163 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2454__B1 _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2057__I0 _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2850__D u0.cmd\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2509__A1 _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2280_ u1.ordering_timer\[2\] _0602_ _0605_ _0619_ _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_42_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2748__A1 _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1995_ net222 _0418_ _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2613__I _0890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1420__A1 u0.cmd\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2616_ _0891_ _0892_ _0893_ _0210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__1971__A2 _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2547_ _0842_ _0192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2478_ _1093_ _0790_ _0791_ _0792_ _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1429_ u1.ordering_complete\[23\] _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_29_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2739__A1 _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output88_I net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2211__I0 _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1714__A2 _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2845__D u0.cmd\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2433__I u1.ordering_timer\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1780_ _1395_ _1396_ _1359_ _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_11_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2202__I0 _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2401_ _1061_ _0720_ _0725_ _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2332_ _0648_ u1.ordering_timer\[9\] _0654_ _0649_ _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2263_ _0603_ _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2194_ _0474_ u1.inverter_select\[7\] _0545_ _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1469__A1 _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1469__B2 u1.ordering_complete\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_36_clock_I clknet_2_0__leaf_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2130__A2 _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2269__I0 u1.ordering_complete\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1641__B2 _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1978_ _0411_ _0412_ _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold13 u0.mem_write_n\[3\] net255 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_0_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold35 u1.inverter_select\[1\] net277 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold24 u1.row_col_select\[8\] net266 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold46 u0.cmd\[3\] net288 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XANTENNA__2970__CLK clknet_leaf_12_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2657__B1 _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output126_I net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1422__I u1.ordering_timer\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2672__A3 _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_15_clock clknet_2_3__leaf_clock clknet_leaf_15_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2360__A2 _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2428__I _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2950_ _0092_ clknet_leaf_4_clock u1.ordering_complete\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2881_ _0015_ clknet_leaf_8_clock u0.mem_write_n\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3259__I clknet_leaf_10_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1901_ u0.cmd\[1\] _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1832_ _0299_ _1160_ _0296_ _0302_ _0015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_31_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2843__CLK clknet_leaf_15_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1763_ _1289_ _1290_ _1379_ _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1694_ _1262_ _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1926__A2 _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2993__CLK clknet_leaf_18_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2315_ _1124_ _0649_ _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3295_ net148 net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2246_ _1057_ _0584_ _0586_ _0587_ _1055_ _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_38_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2338__I _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2103__A2 _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2177_ net218 _0350_ _0452_ _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1614__A1 _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2073__I u0.cmd\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1417__I _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2342__A2 _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2866__CLK clknet_leaf_34_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2333__A2 _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3080_ _0005_ clknet_leaf_12_clock u0.run_state\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1490__C _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2100_ _0491_ _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2031_ _0380_ _0428_ _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1844__A1 _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2933_ _0075_ clknet_leaf_2_clock u1.ccr1\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2864_ net291 clknet_leaf_4_clock control_trigger_sync\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1815_ net19 net37 _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_15_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2795_ _1019_ _0263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3021__CLK clknet_leaf_13_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1746_ _1209_ _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1677_ _1269_ u1.ccr0\[11\] u1.ccr0\[10\] _1268_ _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__3171__CLK clknet_leaf_7_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2269__S _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3278_ net109 net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2068__I u0.cmd\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2229_ _1096_ _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_26_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1835__A1 _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2889__CLK clknet_leaf_3_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_5_clock_I clknet_2_1__leaf_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2531__I _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2179__S _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2315__A2 _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1811__S net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2853__D u0.cmd\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3044__CLK clknet_leaf_1_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2251__A1 _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2441__I u1.ordering_timer\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1600_ u1.ccr1\[1\] _1209_ _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2580_ _1160_ _0858_ _0859_ spi_data_crossing\[27\].data_sync _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_12_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3194__CLK clknet_leaf_30_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1531_ u0.cmd\[29\] _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2597__B _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1462_ u1.ordering_timer\[26\] _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__3272__I net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2089__S _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3201_ _0271_ clknet_leaf_23_clock u1.ccr0\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3132_ net69 net228 spi_data_crossing\[7\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3063_ _0205_ clknet_leaf_6_clock u0.cmd\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2014_ _0431_ _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1520__I _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2490__A1 u1.ordering_complete\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2916_ _0058_ clknet_leaf_26_clock u1.ccr1\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2847_ net288 clknet_leaf_10_clock net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2351__I _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2778_ _1007_ net24 _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1729_ _1177_ _1343_ _1344_ _1345_ _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1505__B1 _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output206_I net206 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3067__CLK clknet_leaf_6_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2481__A1 _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2261__I _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2904__CLK clknet_leaf_36_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2848__D net290 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2436__I _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2472__A1 _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout237_I net238 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2701_ _1295_ _0956_ _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__3267__I net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2632_ _0891_ _0903_ _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput204 net204 row_select_left[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput215 net215 row_select_right[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_2563_ _0846_ _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1514_ _1138_ _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_47_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2494_ u1.ordering_timer\[28\] _0791_ _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1445_ _1057_ _1063_ _1066_ _1069_ _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_3115_ _0249_ clknet_leaf_36_clock u1.timer\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3046_ _0188_ clknet_leaf_1_clock u0.cmd\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2066__I1 u1.ordering_complete\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2927__CLK clknet_leaf_2_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1813__I1 net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3232__CLK clknet_leaf_17_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2367__S _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2693__A1 _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2460__A4 _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1994_ _1271_ _0421_ _0422_ _0059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1420__A2 _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_32_clock_I clknet_2_0__leaf_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2615_ u1.row_sel\[0\] _0875_ _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_47_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2546_ _0388_ _0838_ _0839_ spi_data_crossing\[14\].data_sync _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_47_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2477_ _0780_ _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1428_ _1047_ u1.ordering_complete\[22\] _1049_ u1.ordering_complete\[21\] _1053_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_29_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2076__I u0.cmd\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3029_ _0171_ clknet_leaf_24_clock u1.ordering_timer\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3105__CLK clknet_leaf_31_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2739__A2 _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2675__A1 _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3022__D _0164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2861__D net243 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2400_ _1068_ _0721_ _0724_ _0714_ _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__2202__I1 u1.row_col_select\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2331_ _1109_ _0663_ _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2262_ _0565_ _0600_ _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_2_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3280__I net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2193_ _0548_ _0132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1469__A2 u1.ordering_complete\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1641__A2 _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1977_ _0397_ _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2529_ _0831_ _0185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold14 u0.mem_write_n\[2\] net256 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_29_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold25 u1.inverter_select\[0\] net267 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold36 u1.inverter_select\[8\] net278 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold47 u0.cmd\[5\] net289 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_25_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input32_I la_oenb[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output119_I net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2409__A1 _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2196__I0 _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2856__D net222 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2120__I0 _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2880_ _0014_ clknet_leaf_8_clock u0.mem_write_n\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1900_ _0355_ _0032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2820__A1 net221 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1831_ _0296_ _0302_ _0303_ _0014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_37_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1762_ _1284_ _1288_ _1291_ _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3275__I net106 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1693_ u1.ccr0\[12\] _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_48_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2336__B1 _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2314_ u1.ordering_timer\[6\] u1.ordering_timer\[5\] _0625_ _0628_ _0649_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__and4_1
X_3294_ net146 net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2245_ _1051_ _1053_ _1048_ _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_22_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2176_ _0310_ _0530_ _0538_ _0125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_26_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2111__I0 _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2327__B1 _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1433__I u1.ordering_complete\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_1_clock_I clknet_2_0__leaf_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2264__I _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2802__A1 _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2169__I0 _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2318__B1 _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2030_ _0444_ _0073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3210__D _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2932_ _0074_ clknet_2_0__leaf_clock u1.ccr1\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2863_ net250 clknet_leaf_4_clock control_trigger_sync\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2960__CLK clknet_leaf_20_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1814_ _0292_ _0000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2794_ u1.ccr0\[2\] _0361_ _1017_ _1019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_7_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1745_ _1347_ _1356_ _1361_ _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_15_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1676_ u1.timer\[9\] _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3277_ net108 net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2228_ _1132_ _0568_ _0569_ _1129_ _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_27_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1835__A2 _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2159_ _0393_ _0348_ _0454_ _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_27_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_14_clock clknet_2_3__leaf_clock clknet_leaf_14_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_26_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_29_clock clknet_2_2__leaf_clock clknet_leaf_29_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_6_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2812__I _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2833__CLK clknet_leaf_10_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2983__CLK clknet_leaf_14_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1530_ _1043_ _1152_ _0008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1461_ u1.ordering_complete\[24\] _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_10_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3200_ _0270_ clknet_leaf_31_clock u1.ccr0\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3131_ spi_data_crossing\[6\].A clknet_leaf_0_clock spi_data_crossing\[6\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3062_ _0204_ clknet_leaf_8_clock u0.cmd\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1801__I u1.timer\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2013_ u1.ccr1\[19\] _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_36_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2490__A2 _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2242__A2 _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2915_ _0057_ clknet_leaf_26_clock u1.ccr1\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2846_ u0.cmd\[2\] clknet_leaf_15_clock net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2777_ net6 _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_2_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1728_ u1.timer\[26\] _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1753__A1 _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1659_ _1251_ _1266_ _1276_ _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__2856__CLK clknet_leaf_16_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2079__I u0.cmd\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1505__B2 u1.ordering_complete\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1505__A1 _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_27_clock_I clknet_2_2__leaf_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1808__A2 _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output101_I net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2481__A2 _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1867__B _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3011__CLK clknet_leaf_19_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3161__CLK clknet_leaf_6_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2224__A2 _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2700_ _0945_ _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1983__A1 _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2631_ net216 _0900_ u1.row_sel\[6\] _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_12_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput205 net205 row_select_left[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_2562_ _0844_ _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3283__I net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2879__CLK clknet_leaf_7_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1513_ u1.ordering_timer\[0\] _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2493_ _1082_ u1.ordering_timer\[29\] _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1444_ u1.ordering_timer\[18\] _1067_ _1068_ _1061_ _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_4_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3114_ _0248_ clknet_leaf_36_clock u1.timer\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1531__I u0.cmd\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3045_ _0187_ clknet_leaf_1_clock u0.cmd\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1974__A1 _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2829_ _1038_ _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input62_I spi_data[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3034__CLK clknet_leaf_22_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2151__A1 _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3184__CLK clknet_leaf_33_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2454__A2 _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2859__D net219 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1717__A1 _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1717__B2 _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3278__I net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1993_ _0382_ _0418_ _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1956__A1 _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2614_ u1.row_sel\[0\] _0875_ _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1708__A1 _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3057__CLK clknet_leaf_5_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2545_ _0841_ _0191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2476_ u1.ordering_timer\[27\] _0783_ _1085_ _0784_ _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_1427_ _1048_ _1051_ _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_29_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2133__A1 u0.cmd\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2357__I _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3028_ _0170_ clknet_leaf_24_clock u1.ordering_timer\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1947__A1 _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2372__A1 u1.ordering_complete\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout240 net241 net240 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_8_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2427__A2 u1.ordering_timer\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1938__A1 _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2363__A1 u1.ordering_timer\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2330_ _0654_ _0656_ _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2261_ _0601_ _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2917__CLK clknet_leaf_26_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2192_ _0471_ u1.inverter_select\[6\] _0545_ _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_38_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2126__B _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1976_ u0.cmd\[5\] _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_14_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2354__A1 _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2528_ _0474_ _0826_ _0827_ spi_data_crossing\[7\].data_sync _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold15 u0.mem_write_n\[6\] net257 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold26 u1.col_sel\[0\] net268 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_2459_ _0703_ _0698_ _0775_ _0722_ _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xhold37 u1.u1.impulse_gen\[0\] net279 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_9_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2106__A1 _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold48 u0.cmd\[4\] net290 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XANTENNA_input25_I la_oenb[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2409__A2 _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3222__CLK clknet_leaf_18_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2550__I _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2198__S _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2120__I1 u1.ordering_complete\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1830_ u0.cmd\[26\] _1149_ _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_31_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2584__A1 u0.cmd\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1761_ _1292_ _1369_ _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1692_ _1293_ u1.ccr0\[9\] u1.ccr0\[8\] _1267_ _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2336__A1 u1.ordering_timer\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2313_ u1.ordering_timer\[7\] _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3293_ net144 net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2244_ _1066_ _0585_ _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2175_ _0470_ _0531_ _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_38_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3245__CLK clknet_leaf_8_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2111__I1 u1.ordering_complete\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2370__I u1.ordering_timer\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1959_ u1.ccr1\[0\] _0392_ _0398_ _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2327__A1 _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1915__S _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output131_I net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2802__A2 _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2566__A1 u0.cmd\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2169__I1 u1.col_limit\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2931_ _0073_ clknet_leaf_0_clock u1.ccr1\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2862_ net272 clknet_leaf_5_clock latch_data_sync\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1813_ net18 net1 net36 _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2793_ _1018_ _0262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1744_ _1359_ _1360_ _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2309__A1 u1.ordering_complete\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1675_ _1285_ _1288_ _1291_ _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3276_ net107 net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2227_ _1123_ _1131_ _1126_ _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2158_ _0526_ _0522_ _0527_ _0118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_38_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2089_ _0386_ u1.ordering_complete\[13\] _0456_ _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_41_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1599__A2 u1.ccr1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2548__A1 _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_23_clock_I clknet_2_2__leaf_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2548__B2 spi_data_crossing\[15\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2020__I0 u1.ccr1\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1523__A2 control_trigger vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2087__I0 _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1619__I u1.timer\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1460_ u1.ordering_timer\[24\] _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3090__CLK clknet_leaf_23_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2011__I0 u1.ccr1\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3130_ net68 net228 spi_data_crossing\[6\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2711__A1 _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3061_ _0203_ clknet_leaf_7_clock u0.cmd\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1817__A3 _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2012_ _0433_ _0066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3221__D net282 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2778__A1 _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2914_ _0056_ clknet_leaf_25_clock u1.ccr1\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2845_ u0.cmd\[1\] clknet_leaf_15_clock net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1450__B2 u1.ordering_complete\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2776_ _1006_ net25 _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1727_ u1.ccr0\[26\] _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1658_ u1.ccr1\[8\] _1267_ _1274_ _1275_ _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__1505__A2 u1.ordering_complete\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1589_ _1206_ _1207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3259_ clknet_leaf_10_clock net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_27_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3131__D spi_data_crossing\[6\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1439__I u1.ordering_timer\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1441__A1 _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1441__B2 u1.ordering_complete\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1744__A2 _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2792__I1 _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1902__I _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2950__CLK clknet_leaf_4_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1680__A1 _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2630_ _0891_ _0902_ _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput206 net206 row_select_left[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_2561_ _0851_ _0197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1512_ _1128_ u1.ordering_complete\[3\] _1136_ u1.ordering_complete\[2\] _1137_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
Xclkbuf_leaf_13_clock clknet_2_1__leaf_clock clknet_leaf_13_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_2492_ u1.ordering_complete\[30\] _0792_ _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1443_ u1.ordering_timer\[17\] _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_4_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_28_clock clknet_2_2__leaf_clock clknet_leaf_28_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3113_ _0247_ clknet_leaf_34_clock u1.timer\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2448__B1 _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3044_ _0186_ clknet_leaf_1_clock u0.cmd\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1671__A1 _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1423__B2 u1.ordering_complete\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1974__A2 _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2828_ net13 net31 _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_20_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2759_ _0996_ _0995_ _0997_ _0934_ _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA_input55_I spi_data[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2973__CLK clknet_leaf_11_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2439__B1 _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2553__I _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3036__D _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2846__CLK clknet_leaf_15_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1992_ _0402_ _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_20_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2613_ _0890_ _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3294__I net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2996__CLK clknet_leaf_16_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1708__A2 _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2544_ _0386_ _0838_ _0839_ spi_data_crossing\[13\].data_sync _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2475_ _0783_ _0773_ _0778_ _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1426_ _1049_ u1.ordering_complete\[21\] _1050_ u1.ordering_complete\[20\] _1051_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_25_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2133__A2 _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3027_ _0169_ clknet_leaf_20_clock u1.ordering_timer\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1918__S _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3001__CLK clknet_leaf_17_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2372__A2 _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output161_I net161 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3151__CLK clknet_leaf_5_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout241 net242 net241 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_8_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout230 net232 net230 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_47_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2427__A3 _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2869__CLK clknet_leaf_10_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2260_ _0600_ _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2191_ _0547_ _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1874__A1 _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3024__CLK clknet_leaf_21_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1975_ _1197_ _0403_ _0410_ _0052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2051__A1 _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3174__CLK net240 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2527_ _0830_ _0184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2458_ _0676_ _1116_ _0774_ _0692_ _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_29_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold16 u0.cmd\[22\] net258 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold27 u0.cmd\[17\] net269 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold38 u1.row_col_select\[5\] net280 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_29_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2106__A2 _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold49 control_trigger_sync\[0\] net291 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_2389_ u1.ordering_complete\[16\] _0714_ _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_29_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input18_I la_data_in[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2831__I _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_2_2__f_clock clknet_0_clock clknet_2_2__leaf_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__1447__I u1.ordering_timer\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output86_I net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_18_clock_I clknet_2_3__leaf_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3047__CLK clknet_leaf_1_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2033__A1 _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1760_ _1370_ _1376_ _1368_ _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_11_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3197__CLK clknet_leaf_23_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1691_ _1306_ _1307_ _1308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2336__A2 _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2312_ _0647_ _0152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3292_ net142 net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2243_ _1062_ _1069_ _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2174_ _0537_ _0124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2024__A1 _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1958_ _0397_ _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1889_ u0.cmd\[0\] _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2327__A2 _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2098__I _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1931__S _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2907__CLK clknet_leaf_30_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2810__I0 u1.ccr0\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2318__A2 _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1905__I _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1640__I u1.timer\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2930_ _0072_ clknet_leaf_2_clock u1.ccr1\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2861_ net243 clknet_leaf_5_clock latch_data_sync\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1812_ _0291_ _0002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2792_ u1.ccr0\[1\] _0400_ _1017_ _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_7_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1743_ _1167_ u1.ccr0\[30\] u1.ccr0\[29\] _1168_ _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1765__B1 _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1674_ _1289_ _1290_ _1281_ _1280_ _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2309__A2 _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3275_ net106 net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3212__CLK clknet_leaf_34_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2226_ _1141_ _0567_ _1137_ _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2157_ _0470_ _0516_ _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_27_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2493__A1 _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2088_ _0483_ _0092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2381__I _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3129__D spi_data_crossing\[5\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2020__I1 _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2720__A2 _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2484__A1 _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2087__I1 u1.ordering_complete\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3235__CLK clknet_leaf_7_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2011__I1 _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3060_ _0202_ clknet_leaf_7_clock u0.cmd\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2011_ u1.ccr1\[18\] _0361_ _0432_ _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_35_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3297__I net163 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2913_ _0055_ clknet_leaf_25_clock u1.ccr1\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2844_ u0.cmd\[0\] clknet_leaf_15_clock net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1450__A2 u1.ordering_complete\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2775_ net7 _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1726_ u1.ccr0\[27\] _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1657_ _1247_ _1248_ _1275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_28_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1588_ u1.timer\[0\] _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3258_ clknet_leaf_9_clock net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2376__I _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2209_ _0557_ _0139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3189_ _0259_ clknet_leaf_35_clock net153 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3108__CLK clknet_leaf_31_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1441__A2 u1.ordering_complete\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1729__B1 _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_9_clock clknet_2_1__leaf_clock clknet_leaf_9_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_40_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput207 net207 row_select_left[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_2560_ net218 _0845_ _0847_ spi_data_crossing\[19\].data_sync _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_47_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1511_ u1.ordering_timer\[2\] _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2491_ _1076_ _0709_ _0803_ _0565_ _0175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1442_ u1.ordering_complete\[18\] _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2696__A1 _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3112_ _0246_ clknet_leaf_34_clock u1.timer\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3232__D net266 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3043_ _0185_ clknet_leaf_3_clock u0.cmd\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1671__A2 _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2620__A1 u1.row_sel\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2827_ _1037_ _0277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2758_ _0996_ _0995_ _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1709_ _1324_ _1325_ _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2689_ u1.timer\[7\] u1.timer\[4\] _0941_ _0947_ _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_28_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input48_I spi_data[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2687__A1 _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output204_I net204 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3080__CLK clknet_leaf_12_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1991_ _0420_ _0058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2612_ _0875_ _0889_ _0890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2543_ _0840_ _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2474_ _0789_ _0172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1425_ u1.ordering_timer\[20\] _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_25_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2141__I0 _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3026_ _0168_ clknet_leaf_20_clock u1.ordering_timer\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2940__CLK clknet_leaf_13_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1580__A1 _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2829__I _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1580__B2 u1.timer\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout231 net232 net231 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout220 u0.cmd\[14\] net220 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout242 net72 net242 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_8_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1883__A2 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_12_clock clknet_2_1__leaf_clock clknet_leaf_12_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_42_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1908__I _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_14_clock_I clknet_2_3__leaf_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_27_clock clknet_2_2__leaf_clock clknet_leaf_27_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_13_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2005__S _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2190_ _0468_ u1.inverter_select\[5\] _0545_ _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_38_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2407__C _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2963__CLK clknet_leaf_20_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1974_ _0409_ _0405_ _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2051__A2 _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2526_ _0370_ _0826_ _0827_ spi_data_crossing\[6\].data_sync _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2457_ _0648_ u1.ordering_timer\[9\] _0654_ _0649_ _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_29_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold17 reset_n_sync\[0\] net259 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold28 reset_n net270 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold39 u1.inverter_select\[6\] net281 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_29_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2388_ _0607_ _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3009_ _0151_ clknet_leaf_16_clock u1.ordering_timer\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1617__A2 _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2578__B1 _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2593__A3 _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2836__CLK clknet_leaf_10_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2986__CLK clknet_leaf_16_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2033__A2 _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1638__I u1.timer\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1792__A1 _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1690_ _1256_ u1.ccr0\[15\] u1.ccr0\[14\] _1257_ _1307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2311_ u1.ordering_timer\[6\] _0627_ _0635_ _0646_ _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1544__A1 _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3291_ net140 net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2242_ _0583_ _1058_ _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2173_ _0468_ u1.col_limit\[5\] _0529_ _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1480__B1 u1.ordering_timer\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2024__A2 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3141__CLK clknet_leaf_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1957_ _0396_ _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1888_ _0331_ _0344_ _0031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1783__A1 _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2859__CLK clknet_leaf_16_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2509_ _1042_ u0.latch_cmd _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input30_I la_oenb[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1838__A2 _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2810__I1 _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3014__CLK clknet_leaf_21_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1921__I _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3164__CLK net239 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2860_ net249 clknet_leaf_9_clock net192 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1811_ net17 net2 net35 _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_19_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2791_ _1011_ _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1742_ u1.timer\[29\] _1357_ _1358_ u1.timer\[28\] _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_15_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1673_ u1.ccr0\[7\] _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3274_ net105 net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2225_ _1135_ _1140_ _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2156_ u1.row_limit\[6\] _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2087_ _0447_ u1.ordering_complete\[12\] _0456_ _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2989_ _0131_ clknet_leaf_18_clock u1.inverter_select\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1756__A1 _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3145__D spi_data_crossing\[13\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3037__CLK clknet_leaf_3_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1741__I u1.ccr0\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3187__CLK clknet_leaf_33_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1692__B1 u1.ccr0\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2572__I _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1444__B1 _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1995__A1 net222 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2010_ _0431_ _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2475__A2 _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2912_ _0054_ clknet_leaf_24_clock u1.ccr1\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2843_ u1.col_sel\[5\] clknet_leaf_15_clock net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2774_ _1005_ net26 _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1738__A1 _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1725_ _1323_ _1326_ _1341_ _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1656_ u1.ccr1\[10\] _1268_ _1270_ _1273_ _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1587_ u1.ccr1\[2\] _1204_ _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2163__A1 _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1910__A1 _1320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3257_ clknet_leaf_9_clock net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2208_ _0364_ u1.row_col_select\[3\] _0553_ _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3188_ _0258_ clknet_leaf_33_clock net155 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2139_ _0347_ _0348_ _0454_ _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_26_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1426__B1 _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2154__A1 _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2457__A2 u1.ordering_timer\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2235__C _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1968__A1 _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3202__CLK clknet_leaf_23_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput208 net208 row_select_left[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__2251__B _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1510_ u1.ordering_timer\[0\] _1133_ u1.ordering_timer\[1\] _1134_ _1135_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_2490_ u1.ordering_complete\[29\] _0720_ _0709_ _0802_ _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1441_ _1064_ u1.ordering_complete\[19\] _1065_ u1.ordering_complete\[18\] _1066_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_4_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2477__I _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3111_ _0245_ clknet_leaf_34_clock u1.timer\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2696__A2 _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3042_ _0184_ clknet_leaf_3_clock u0.cmd\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2448__A2 _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2826_ net4 net22 _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_20_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2757_ u1.timer\[29\] _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2688_ _0946_ _0948_ _0949_ _0226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1708_ _1318_ _1319_ _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1639_ u1.timer\[14\] _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2136__A1 _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2687__A2 _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3309_ net206 net212 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2439__A2 _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3225__CLK clknet_leaf_17_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2297__I _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2678__A2 _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_10_clock_I clknet_2_1__leaf_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1990_ u1.ccr1\[10\] _0380_ _0402_ _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_18_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2602__A2 _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout228_I net229 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2611_ _0886_ _0887_ _0888_ _0329_ _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_9_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2542_ _0447_ _0838_ _0839_ spi_data_crossing\[12\].data_sync _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_5_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2118__A1 u0.cmd\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2473_ _0783_ _0716_ _0761_ _0788_ _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1424_ u1.ordering_timer\[21\] _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2892__CLK clknet_leaf_2_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3248__CLK clknet_leaf_9_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3025_ _0167_ clknet_leaf_20_clock u1.ordering_timer\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_8_clock clknet_2_1__leaf_clock clknet_leaf_8_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_30_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2809_ _1027_ _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input60_I spi_data[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2111__S _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2109__A1 _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout221 u0.cmd\[13\] net221 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout232 net233 net232 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_47_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2348__A1 u1.ordering_complete\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1924__I u0.cmd\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1973_ u0.cmd\[4\] _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3238__D u0.cmd\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2339__A1 u1.ordering_timer\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2525_ _0829_ _0183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_29_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2456_ u1.ordering_timer\[25\] _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold29 u1.row_sel\[4\] net271 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold18 u1.row_col_select\[9\] net260 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XANTENNA__3070__CLK clknet_leaf_9_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2387_ _1059_ _0712_ _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_25_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3008_ _0150_ clknet_leaf_14_clock u1.ordering_timer\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1928__I1 _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3093__CLK clknet_leaf_26_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2310_ _0643_ _0644_ _0645_ _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3290_ net157 net156 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2741__A1 _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2241_ u1.ordering_timer\[19\] _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2172_ _0536_ _0123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2930__CLK clknet_leaf_2_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1480__B2 _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1956_ _0393_ _0395_ _0351_ _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1887_ u1.col_sel\[6\] _0343_ _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2732__A1 _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2508_ _0817_ _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_11_clock clknet_2_1__leaf_clock clknet_leaf_11_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_2439_ _0753_ _0754_ _0733_ _0758_ _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_29_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input23_I la_oenb[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2395__I _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_26_clock clknet_2_2__leaf_clock clknet_leaf_26_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_16_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2799__A1 _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2953__CLK clknet_leaf_3_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1810_ _0290_ _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_19_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2790_ _1010_ _1014_ _1016_ _0261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_8_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1741_ u1.ccr0\[28\] _1358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1672_ u1.timer\[7\] _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1517__A2 u1.ordering_complete\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2714__A1 _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3273_ net104 net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2224_ _1070_ _1095_ _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2155_ _0524_ _0522_ _0525_ _0117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_6_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2086_ _1104_ _0457_ _0482_ _0091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_19_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2988_ _0130_ clknet_leaf_18_clock u1.inverter_select\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2402__B1 _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1939_ _1343_ _0379_ _0383_ _0043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2611__C _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2005__I0 u1.ccr1\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2976__CLK clknet_leaf_11_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2705__A1 _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1692__A1 _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1692__B2 _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1444__B2 _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1444__A1 u1.ordering_timer\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1995__A2 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3131__CLK clknet_leaf_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2475__A3 _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2849__CLK clknet_leaf_16_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2911_ _0053_ clknet_leaf_24_clock u1.ccr1\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2842_ net294 clknet_leaf_15_clock net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2773_ net8 _1005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2204__S _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2999__CLK clknet_leaf_18_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1738__A2 u1.ccr0\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1724_ _1333_ _1334_ _1335_ _1340_ _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_1655_ _1271_ _1272_ u1.ccr1\[10\] _1268_ _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1586_ _1203_ _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2163__A2 _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3256_ clknet_leaf_9_clock net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1910__A2 _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2207_ _0556_ _0138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3187_ _0257_ clknet_leaf_33_clock net157 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2138_ _1073_ _0492_ _0514_ _0111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2069_ _0470_ _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1426__B2 u1.ordering_complete\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3004__CLK clknet_leaf_13_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1729__A2 _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2154__A2 _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold1_I latch_data vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2457__A3 _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2583__I _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1968__A2 _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2217__I0 _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1927__I u0.cmd\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2393__A2 _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput209 net209 row_select_left[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_1440_ u1.ordering_timer\[18\] _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1662__I _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3110_ _0244_ clknet_leaf_33_clock u1.timer\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3041_ _0183_ clknet_leaf_4_clock u0.cmd\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1656__A1 u1.ccr1\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2605__B1 u1.row_limit\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3027__CLK clknet_leaf_20_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2208__I0 _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2825_ _1304_ _1015_ _1036_ _0276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3177__CLK clknet_leaf_7_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2756_ _0982_ _0994_ _0995_ _0248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1707_ _1321_ _1320_ _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2687_ _1283_ _0942_ _1280_ _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1638_ u1.timer\[15\] _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1592__B1 u1.ccr1\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2136__A2 _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1569_ _1170_ _1175_ _1182_ _1186_ _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_3308_ net205 net211 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1505__C _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3239_ u0.cmd\[21\] clknet_leaf_7_clock net167 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1583__B1 _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1431__B _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2610_ u1.row_sel\[6\] _0526_ _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2366__A2 _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2541_ _0820_ _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2472_ _0711_ _0786_ _0787_ _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1574__B1 u1.ccr1\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1423_ _1046_ u1.ordering_complete\[23\] _1047_ u1.ordering_complete\[22\] _1048_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__2118__A2 _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3024_ _0166_ clknet_leaf_21_clock u1.ordering_timer\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2054__A1 _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2808_ u1.ccr0\[8\] _0375_ _1013_ _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2739_ _0286_ _0981_ _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_input53_I spi_data[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2109__A2 _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout222 u0.cmd\[12\] net222 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout233 net242 net233 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_28_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2293__A1 u1.ordering_complete\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2045__A1 u0.cmd\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2348__A2 _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1556__B1 u1.ccr1\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1940__I _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2284__A1 _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout240_I net241 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1972_ _1213_ _0403_ _0408_ _0051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_18_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2339__A2 _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2524_ _0368_ _0826_ _0827_ spi_data_crossing\[5\].data_sync _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3215__CLK clknet_leaf_17_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2455_ _0772_ _0170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold19 u1.inverter_select\[5\] net261 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_2386_ _0703_ _0698_ _0694_ _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_25_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1850__I u1.col_sel\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3007_ _0149_ clknet_leaf_12_clock u1.ordering_timer\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_25_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2290__A4 u1.ordering_timer\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2578__A2 _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2122__S _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2792__S _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2882__CLK clknet_leaf_8_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3238__CLK clknet_leaf_7_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1792__A3 _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2240_ _1202_ _1277_ _0579_ _0581_ _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_2171_ _0466_ u1.col_limit\[4\] _0529_ _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1670__I u1.timer\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_7_clock clknet_2_1__leaf_clock clknet_leaf_7_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_4_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2257__A1 _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1480__A2 _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1955_ _0394_ _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_21_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1886_ u1.col_sel\[5\] _0340_ _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2507_ _0816_ _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2438_ _0734_ _0755_ _0757_ _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_9_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2369_ _0697_ _0159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_45_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1838__A4 _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2248__A1 _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input16_I la_data_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2799__A2 _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3300__I net166 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2420__A1 u1.ordering_complete\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2723__A2 u1.timer\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2487__A1 u1.ordering_timer\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2239__A1 _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3060__CLK clknet_leaf_7_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1740_ u1.ccr0\[29\] _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_8_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1671_ _1283_ _1282_ _1286_ _1287_ _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2714__A2 _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3272_ net103 net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input8_I la_data_in[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2223_ _1402_ _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2478__A1 _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2154_ _0411_ _0516_ _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2085_ net223 _0480_ _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_19_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2650__A1 _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2987_ _0129_ clknet_leaf_18_clock u1.inverter_select\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2402__A1 _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1938_ _0382_ _0371_ _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1869_ u0.timer_enable _0309_ _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1575__I u1.timer\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2005__I1 _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1692__A2 u1.ccr0\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3083__CLK clknet_leaf_4_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1485__I u1.ordering_complete\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2920__CLK clknet_leaf_28_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold24_I u1.row_col_select\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2632__A1 _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2910_ _0052_ clknet_leaf_24_clock u1.ccr1\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_10_clock clknet_2_1__leaf_clock clknet_leaf_10_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_2841_ u1.col_sel\[3\] clknet_leaf_15_clock net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2772_ _1004_ net27 _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1723_ _1336_ _1337_ _1338_ _1339_ _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xclkbuf_leaf_25_clock clknet_2_2__leaf_clock clknet_leaf_25_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1654_ u1.timer\[11\] _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2699__A1 _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1585_ u1.timer\[2\] _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3255_ clknet_leaf_9_clock net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2206_ _0461_ u1.row_col_select\[2\] _0553_ _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2171__I0 _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3186_ _0256_ clknet_leaf_33_clock net140 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1674__A2 _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2137_ u0.cmd\[15\] _0509_ _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_35_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2068_ u0.cmd\[6\] _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1426__A2 u1.ordering_complete\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2943__CLK clknet_leaf_14_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3172__D net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2311__B1 _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2457__A4 _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2614__A1 u1.row_sel\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2217__I1 u1.row_col_select\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1943__I net221 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2040__S _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3040_ _0182_ clknet_leaf_4_clock u0.cmd\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1656__A2 _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2966__CLK clknet_leaf_3_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2215__S _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2824_ net219 _1017_ _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2755_ _1413_ _0993_ _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2014__I _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2686_ _0942_ _0947_ _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1706_ _1318_ _1319_ _1320_ _1322_ _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_1637_ _1252_ u1.timer\[15\] _1253_ _1254_ _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_28_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3307_ net204 net210 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1568_ _1183_ _1184_ _1185_ _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1499_ u1.ordering_timer\[7\] _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3238_ u0.cmd\[20\] clknet_leaf_7_clock net166 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3169_ spi_data_crossing\[25\].A clknet_leaf_7_clock spi_data_crossing\[25\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2684__I _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3121__CLK clknet_leaf_35_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1583__A1 _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1583__B2 _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2839__CLK clknet_leaf_10_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1886__A2 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2989__CLK clknet_leaf_18_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2540_ _0817_ _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2471_ u1.ordering_complete\[26\] _0756_ _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1574__A1 u1.ccr1\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1422_ u1.ordering_timer\[22\] _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_25_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3023_ _0165_ clknet_leaf_21_clock u1.ordering_timer\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2826__A1 net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2009__I _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2054__A2 _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2807_ _1290_ _1025_ _1026_ _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2738_ _0286_ _0981_ _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1565__A1 u1.ccr1\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2669_ _1364_ _1208_ _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_input46_I spi_data[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout223 u0.cmd\[11\] net223 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout234 net236 net234 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_41_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3303__I net169 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2293__A2 _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1556__B2 _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3017__CLK clknet_leaf_13_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3167__CLK clknet_leaf_7_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout233_I net242 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1971_ _0407_ _0405_ _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2523_ _0828_ _0182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2454_ _0768_ _0754_ _0761_ _0771_ _0772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2385_ _0608_ _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput1 io_control_trigger_in net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_37_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3006_ _0148_ clknet_leaf_12_clock u1.ordering_timer\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_25_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1578__I u1.ccr1\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1786__A1 _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3180__D net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1474__B1 u1.ordering_timer\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1488__I u1.ordering_complete\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2170_ _0535_ _0122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2662__C1 _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1954_ u0.cmd\[17\] _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1768__A1 _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1885_ _0331_ _0342_ _0030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_31_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2506_ _0815_ u0.latch_cmd _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2437_ u1.ordering_complete\[22\] _0756_ _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2368_ u1.ordering_timer\[13\] _0682_ _0691_ _0696_ _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2496__A2 _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2299_ u1.ordering_timer\[5\] _0625_ _0628_ _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_38_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2248__A2 _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2420__A2 _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2723__A3 _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput190 net190 mem_write_n[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2487__A2 _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1695__B1 _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_21_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3205__CLK clknet_leaf_23_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1946__I net220 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1670_ u1.timer\[4\] _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3085__D _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2175__A1 _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1922__A1 _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3271_ net102 net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2222_ _0564_ _0145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2478__A2 _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2153_ u1.row_limit\[5\] _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2084_ _1113_ _0457_ _0481_ _0090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_35_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1438__B1 _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2650__A2 _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2986_ _0128_ clknet_leaf_16_clock u1.inverter_select\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2402__A2 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1937_ net223 _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1868_ _0330_ _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput70 spi_data[8] net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_1799_ _1318_ _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1913__A1 _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2872__CLK clknet_leaf_14_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3228__CLK clknet_leaf_17_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2641__A2 _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_6_clock clknet_2_1__leaf_clock clknet_leaf_6_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_10_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2157__A1 _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2038__S _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2840_ net225 clknet_leaf_15_clock net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2771_ net9 _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_8_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1722_ _1237_ u1.ccr0\[16\] _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1653_ u1.ccr1\[11\] _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1584_ _1192_ _1195_ _1198_ _1201_ _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__2895__CLK clknet_leaf_3_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3254_ clknet_leaf_9_clock net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2205_ _0555_ _0137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2171__I1 u1.col_limit\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3185_ _0255_ clknet_leaf_33_clock net142 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2136_ _1078_ _0492_ _0513_ _0110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2067_ _0469_ _0085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2623__A2 _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1586__I _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2969_ _0111_ clknet_leaf_22_clock u1.ordering_complete\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2387__A1 _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3306__I net192 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2210__I _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2311__A1 u1.ordering_timer\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3050__CLK clknet_leaf_1_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2366__B _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2614__A2 _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2378__A1 _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2823_ _1305_ _1015_ _1035_ _0275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2754_ _1413_ _0993_ _0994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1705_ _1321_ _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2685_ u1.timer\[6\] u1.timer\[5\] _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_28_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1636_ u1.timer\[14\] _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1592__A2 u1.ccr1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3073__CLK clknet_leaf_10_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1567_ u1.ccr1\[31\] _1171_ _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3306_ net192 net193 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1498_ _1121_ u1.ordering_complete\[5\] _1122_ u1.ordering_complete\[4\] _1123_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3237_ net218 clknet_leaf_7_clock net165 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3168_ net57 net237 spi_data_crossing\[25\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2119_ _1054_ _0502_ _0503_ _0103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_15_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3099_ _0233_ clknet_leaf_29_clock u1.timer\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2910__CLK clknet_leaf_24_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2080__I0 _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2141__S _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2780__A1 _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1583__A2 u1.timer\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3183__D _0253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2532__A1 _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2532__B2 spi_data_crossing\[8\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_24_clock clknet_2_2__leaf_clock clknet_leaf_24_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_46_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2071__I0 _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1954__I u0.cmd\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3096__CLK clknet_leaf_27_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2470_ _1087_ _0785_ _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1421_ u1.ordering_timer\[23\] _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_1_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2933__CLK clknet_leaf_2_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2785__I _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3022_ _0164_ clknet_leaf_30_clock u1.ordering_timer\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2806_ _0373_ _1021_ _1026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2737_ _0933_ _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2668_ _1206_ _0935_ _0220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1619_ u1.timer\[16\] _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2599_ u1.row_sel\[3\] _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2514__B2 spi_data_crossing\[1\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2514__A1 _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout235 net236 net235 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_8_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout224 u0.cmd\[10\] net224 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input39_I la_oenb[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2753__A1 _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2956__CLK clknet_leaf_3_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1492__A1 _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1492__B2 u1.ordering_complete\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1949__I net219 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1970_ u0.cmd\[3\] _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2522_ _0366_ _0826_ _0827_ spi_data_crossing\[4\].data_sync _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2744__A1 u1.timer\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2453_ _0734_ _0769_ _0770_ _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2384_ _0709_ _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput2 io_latch_data_in net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3005_ _0147_ clknet_leaf_12_clock u1.ordering_timer\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3111__CLK clknet_leaf_34_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1786__A2 _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1594__I u0.timer_enable vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2979__CLK clknet_leaf_14_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1474__B2 _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1474__A1 _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2726__A1 _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold47_I u0.cmd\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1465__A1 _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1953_ u0.cmd\[16\] _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1884_ _0311_ _0340_ _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_30_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2717__A1 _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2505_ _1041_ _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2436_ _0596_ _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2367_ u1.ordering_complete\[13\] _0695_ _0609_ _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_29_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2298_ _0634_ _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3007__CLK clknet_leaf_12_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3309__I net206 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2708__A1 _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3157__CLK clknet_leaf_5_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput180 net180 mem_address_right[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput191 net191 mem_write_n[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_48_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1695__B2 _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1998__A2 _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2644__B1 _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2175__A2 _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3270_ net95 net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2221_ _0478_ u1.row_col_select\[9\] _0552_ _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2152_ _0521_ _0522_ _0523_ _0116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_26_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2083_ net224 _0480_ _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_35_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1438__A1 u1.ordering_timer\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1438__B2 _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2985_ _0127_ clknet_leaf_16_clock u1.inverter_select\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1936_ _1344_ _0379_ _0381_ _0042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1867_ _0309_ _0328_ _0329_ _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinput60 spi_data[28] net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput71 spi_data[9] net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_1798_ _1412_ _1414_ _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2166__A2 _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1913__A2 _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2419_ _1050_ _0736_ _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_40_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input21_I la_data_in[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1677__B2 _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1677__A1 _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output108_I net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2652__B _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3186__D _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2157__A2 _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1668__B2 _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1668__A1 _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1450__C _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2093__A1 net219 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1840__A1 _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1957__I _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2770_ _1003_ net28 _0254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1721_ _1224_ u1.ccr0\[20\] _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1652_ u1.ccr1\[11\] _1269_ _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2788__I _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1583_ _1199_ u1.timer\[7\] _1200_ _1188_ _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3253_ net244 clknet_leaf_9_clock net191 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2204_ _0357_ u1.row_col_select\[1\] _0553_ _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3184_ _0254_ clknet_leaf_33_clock net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2135_ u0.cmd\[14\] _0509_ _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_26_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2066_ _0468_ u1.ordering_complete\[5\] _0462_ _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_19_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2084__A1 _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2028__I _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2968_ _0110_ clknet_leaf_22_clock u1.ordering_complete\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1919_ _0369_ _0037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2899_ _0041_ clknet_leaf_36_clock u1.ccr0\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2139__A2 _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input69_I spi_data[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2311__A2 _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2822_ net220 _1017_ _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2862__CLK clknet_leaf_5_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2753_ _0983_ _0992_ _0993_ _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1704_ u1.timer\[18\] _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2684_ _0945_ _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3218__CLK clknet_leaf_17_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1635_ u1.ccr1\[14\] _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1566_ u1.ccr1\[28\] _1173_ u1.ccr1\[24\] _1165_ _1184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3305_ net171 net181 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1497_ u1.ordering_timer\[4\] _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3236_ u0.cmd\[18\] clknet_leaf_7_clock net164 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3167_ spi_data_crossing\[24\].A clknet_leaf_7_clock spi_data_crossing\[24\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_5_clock clknet_2_1__leaf_clock clknet_leaf_5_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_2118_ u0.cmd\[7\] _0495_ _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3098_ _0232_ clknet_leaf_27_clock u1.timer\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2049_ _0456_ _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_8_clock_I clknet_2_1__leaf_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2080__I1 _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2885__CLK clknet_leaf_8_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2071__I1 u1.ordering_complete\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1420_ u0.cmd\[26\] _1044_ _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1970__I u0.cmd\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1731__B1 u1.ccr0\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3021_ _0163_ clknet_leaf_13_clock u1.ordering_timer\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2805_ _1012_ _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3040__CLK clknet_leaf_4_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2736_ _1233_ _0980_ _0981_ _0982_ _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2667_ _0934_ _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1618_ u1.timer\[17\] _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2598_ net217 _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3190__CLK clknet_leaf_35_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout225 u1.col_sel\[2\] net225 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_1549_ u1.timer\[30\] _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
Xfanout236 net241 net236 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_45_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3219_ net261 clknet_leaf_17_clock net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1713__B1 _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1492__A2 u1.ordering_complete\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3063__CLK clknet_leaf_6_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1965__I _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout219_I u0.cmd\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2521_ _0820_ _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2900__CLK clknet_leaf_34_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2452_ u1.ordering_complete\[24\] _0756_ _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2383_ _0601_ _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_25_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3004_ _0146_ clknet_leaf_13_clock u1.ordering_timer\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput3 io_reset_n_in net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_36_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2680__A1 _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2480__B _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2719_ _0968_ _0969_ _0971_ _0235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
Xclkbuf_leaf_23_clock clknet_2_2__leaf_clock clknet_leaf_23_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_47_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input51_I spi_data[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2147__S _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1474__A2 _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3086__CLK clknet_leaf_29_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3189__D _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1785__I _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2026__I1 _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2923__CLK clknet_leaf_2_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2057__S _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2662__A1 u1.ccr1\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1952_ u0.cmd\[0\] _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1883_ _0330_ _0340_ _0341_ _0029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_30_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2717__A2 _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_35_clock_I clknet_2_0__leaf_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2504_ _0810_ _0709_ _0814_ _0177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2435_ _1047_ _0749_ _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_9_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2350__B1 _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2366_ _1101_ _0685_ _0694_ _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2297_ _0603_ _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2946__CLK clknet_leaf_19_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2405__A1 _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1613__C1 u1.ccr1\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2708__A2 _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2430__S _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput170 net170 mem_address_left[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput181 net181 mem_address_right[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput192 net192 output_active_left vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2192__I0 _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2644__A1 _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3101__CLK clknet_leaf_28_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2580__B1 _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3251__CLK clknet_leaf_9_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2220_ _0563_ _0144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2183__I0 _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2151_ _0409_ _0522_ _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_26_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2082_ _0455_ _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1438__A2 _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2969__CLK clknet_leaf_22_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2984_ _0126_ clknet_leaf_18_clock u1.inverter_select\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2742__C _0982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1935_ _0380_ _0371_ _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1866_ _1402_ _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput61 spi_data[29] net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput50 spi_data[19] net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput72 spi_data_clock net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_1797_ _1351_ u1.timer\[30\] u1.timer\[29\] _1413_ _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_1_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2418_ _0740_ _0165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2349_ _0670_ _0678_ _0679_ _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input14_I la_data_in[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2626__A1 net217 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2617__A1 _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1720_ _1233_ u1.ccr0\[21\] _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1973__I u0.cmd\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1651_ u1.timer\[11\] _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_7_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1582_ u1.ccr1\[6\] _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3252_ net246 clknet_leaf_9_clock net190 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2203_ _0554_ _0136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2305__B1 _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input6_I la_data_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3183_ _0253_ clknet_leaf_28_clock net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1659__A2 _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2134_ _1079_ _0502_ _0512_ _0109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_27_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2608__B2 net217 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2065_ _0411_ _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_19_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2084__A2 _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3147__CLK clknet_leaf_1_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2967_ _0109_ clknet_leaf_23_clock u1.ordering_complete\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2898_ _0040_ clknet_leaf_0_clock u1.ccr0\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1918_ u1.ccr0\[21\] _0368_ _0354_ _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1849_ _0311_ u1.col_limit\[5\] _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_33_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2147__I0 _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2647__C _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_4_clock_I clknet_2_1__leaf_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1510__B2 _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2821_ _1301_ _1015_ _1034_ _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2752_ _1394_ _1345_ _1411_ _0988_ _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__1577__B2 _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1703_ u1.ccr0\[18\] _1320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1577__A1 u1.ccr1\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2683_ _0933_ _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1634_ u1.ccr1\[15\] _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_28_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1565_ u1.ccr1\[25\] _1163_ _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3304_ net170 net180 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3235_ net269 clknet_leaf_7_clock net163 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1496_ u1.ordering_timer\[5\] _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3166_ net56 net237 spi_data_crossing\[24\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1501__A1 _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1501__B2 u1.ordering_complete\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2117_ _0489_ _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3097_ _0231_ clknet_leaf_26_clock u1.timer\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2048_ _0455_ _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_11_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output168_I net168 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2658__B _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3020_ _0162_ clknet_leaf_13_clock u1.ordering_timer\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1899__S _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2804_ _1281_ _1014_ _1024_ _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2750__C _0982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2735_ _0945_ _0982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2666_ _0933_ _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1617_ u1.ccr1\[20\] _1224_ _1232_ _1234_ _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_2597_ _0309_ _0874_ _1212_ _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xfanout226 u1.col_sel\[0\] net226 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout237 net238 net237 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__2478__B _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1548_ _1165_ _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__1722__A1 _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1479_ u1.ordering_complete\[11\] _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_3218_ net262 clknet_leaf_17_clock net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2278__A2 _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3149_ spi_data_crossing\[15\].A clknet_leaf_1_clock spi_data_crossing\[15\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2753__A3 _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2852__CLK clknet_leaf_16_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3208__CLK clknet_leaf_35_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1795__A4 u1.timer\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2744__A3 _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2520_ _0817_ _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_4_clock clknet_2_1__leaf_clock clknet_leaf_4_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_2451_ _0768_ _0764_ _0769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_29_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2382_ _1059_ _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_25_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3003_ _0145_ clknet_leaf_18_clock u1.row_col_select\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput4 la_data_in[0] net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_37_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_31_clock_I clknet_2_0__leaf_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2680__A2 _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2718_ _0970_ _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1891__I u0.cmd\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2649_ _1277_ _0916_ _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2875__CLK clknet_leaf_4_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input44_I spi_data[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2726__A3 u1.timer\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3030__CLK clknet_leaf_24_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2662__A2 _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3180__CLK net240 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1976__I u0.cmd\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2414__A2 _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1951_ _1352_ _0362_ _0391_ _0047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1882_ u1.col_sel\[4\] _0338_ _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_31_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2503_ _0604_ _0813_ _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2898__CLK clknet_leaf_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1925__A1 _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2600__I u1.row_sel\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2434_ _0601_ _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2365_ _0693_ _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2350__A1 _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2296_ _0633_ _0150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2102__A1 _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2405__A2 _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput160 net160 io_update_cycle_complete_oeb vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput182 net182 mem_write_n[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput171 net171 mem_address_left[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput193 net193 output_active_right vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__3053__CLK clknet_leaf_5_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2341__A1 _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2644__A2 _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2580__A1 _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2150_ _0515_ _0522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2081_ _0479_ _0089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_22_clock clknet_2_2__leaf_clock clknet_leaf_22_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_37_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2983_ _0125_ clknet_leaf_14_clock u1.col_limit\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1934_ net224 _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_37_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1865_ u1.col_sel\[6\] _0310_ _0327_ _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xinput40 spi_data[0] net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput51 spi_data[1] net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput62 spi_data[2] net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_1796_ u1.timer\[28\] _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3076__CLK clknet_leaf_5_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2417_ _0583_ _0719_ _0733_ _0739_ _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_44_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2348_ u1.ordering_complete\[11\] _0658_ _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_45_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2279_ _0613_ _0617_ _0618_ _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_26_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2913__CLK clknet_leaf_25_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2505__I _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_0_clock_I clknet_2_0__leaf_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2314__A1 u1.ordering_timer\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1840__A3 _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3099__CLK clknet_leaf_29_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1650_ u1.timer\[10\] _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1581_ u1.ccr1\[7\] _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2150__I _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3251_ net245 clknet_leaf_9_clock net189 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2936__CLK clknet_leaf_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2202_ _0346_ u1.row_col_select\[0\] _0553_ _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3182_ _0252_ clknet_leaf_32_clock net148 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2133_ u0.cmd\[13\] _0509_ _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1903__I1 _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2608__A2 net216 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2064_ _0467_ _0084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2966_ _0108_ clknet_leaf_3_clock u1.ordering_complete\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1917_ u0.cmd\[5\] _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2897_ _0039_ clknet_leaf_2_clock u1.ccr0\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1848_ u1.col_sel\[5\] _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_2_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1779_ _1350_ _1347_ _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2544__A1 _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2663__C _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3241__CLK clknet_leaf_7_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2171__S _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2959__CLK clknet_leaf_20_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1510__A2 _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2820_ net221 _1029_ _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2074__I0 _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2751_ _1410_ _0990_ _1394_ _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_9_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2774__A1 _1005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2682_ _0935_ _0944_ _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1702_ u1.ccr0\[19\] _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1577__A2 _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1633_ _1247_ _1248_ _1249_ _1250_ _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2526__A1 _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1564_ _1176_ _1177_ _1179_ _1181_ _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__2526__B2 spi_data_crossing\[6\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3303_ net169 net179 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1495_ _1108_ _1115_ _1119_ _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_28_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3234_ u0.cmd\[16\] clknet_leaf_7_clock net162 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3114__CLK clknet_leaf_36_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1501__A2 u1.ordering_complete\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3165_ spi_data_crossing\[23\].A clknet_leaf_6_clock spi_data_crossing\[23\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2116_ _0501_ _0102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3096_ _0230_ clknet_leaf_27_clock u1.timer\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2047_ _0452_ _0454_ _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2055__I _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2949_ _0091_ clknet_leaf_12_clock u1.ordering_complete\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_26_clock_I clknet_2_2__leaf_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2756__A1 _0982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3137__CLK clknet_leaf_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1731__A2 u1.ccr0\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1495__A1 _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1798__A2 _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2803_ _0470_ _1021_ _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2603__I u1.row_sel\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2734_ u1.timer\[21\] u1.timer\[20\] _0281_ _0976_ _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_2665_ _1279_ _0932_ _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2596_ _0320_ _0872_ _0873_ _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1616_ u1.ccr1\[21\] _1233_ u1.ccr1\[20\] _1223_ _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_5_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout216 u1.row_sel\[5\] net216 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout238 net239 net238 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__2478__C _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout227 net229 net227 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_1547_ u1.timer\[24\] _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1478_ u1.ordering_timer\[12\] _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3217_ net253 clknet_leaf_16_clock net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3148_ net46 net234 spi_data_crossing\[15\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1889__I u0.cmd\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3079_ _0004_ clknet_leaf_12_clock u0.run_state\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2738__A1 _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2513__I _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1713__A2 _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1477__A1 _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1477__B2 u1.ordering_complete\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1799__I _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2029__I0 u1.ccr1\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2744__A4 _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2450_ _1085_ _0768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3254__I clknet_leaf_9_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2381_ _0707_ _0161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_49_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3002_ _0144_ clknet_leaf_18_clock u1.row_col_select\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput5 la_data_in[10] net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_37_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2417__B1 _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2717_ _1303_ _0966_ _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2648_ _0911_ _0913_ _0915_ _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2489__B _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2579_ _0862_ _0204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input37_I la_oenb[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2508__I _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2726__A4 _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1950_ _0390_ _0384_ _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1881_ u1.col_sel\[4\] _0338_ _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_41_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1622__A1 u1.ccr1\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout224_I u0.cmd\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1992__I _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2502_ u1.ordering_complete\[31\] _0812_ _0780_ _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2433_ u1.ordering_timer\[22\] _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2364_ _0676_ _1116_ _0665_ _0692_ _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_29_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1689__A1 _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1689__B2 _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2350__A2 _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2295_ _0625_ _0627_ _0605_ _0632_ _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_42_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2638__B1 u1.ccr1\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2102__A2 _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1861__B2 u1.col_limit\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1613__A1 u1.ccr1\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2842__CLK clknet_leaf_15_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput150 net150 io_driver_io_oeb[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput161 net161 io_update_cycle_complete_out vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput183 net183 mem_write_n[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput194 net194 row_col_select[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput172 net172 mem_address_right[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__2992__CLK clknet_leaf_18_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_3_clock clknet_2_1__leaf_clock clknet_leaf_3_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_16_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1852__B2 u1.col_limit\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1604__A1 _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold45_I u1.row_col_select\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2580__A2 _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2332__A2 u1.ordering_timer\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2080_ _0478_ _1110_ _0472_ _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_47_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1987__I _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2982_ _0124_ clknet_leaf_16_clock u1.col_limit\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2865__CLK clknet_leaf_33_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1933_ _0359_ _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1864_ _0312_ _0325_ _0326_ _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xinput30 la_oenb[17] net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput63 spi_data[30] net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput52 spi_data[20] net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_1795_ _1394_ _1410_ _1411_ u1.timer\[24\] _1412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
Xinput41 spi_data[10] net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_2416_ _0734_ _0737_ _0738_ _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2347_ _0676_ _0677_ _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_38_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2278_ u1.ordering_complete\[2\] _0597_ _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_29_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1834__A1 _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1897__I _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3020__CLK clknet_leaf_13_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2521__I _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2169__S _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2888__CLK clknet_leaf_3_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1580_ _1196_ _1190_ _1197_ u1.timer\[4\] _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3250_ net257 clknet_leaf_8_clock net188 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3262__I clknet_leaf_10_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2201_ _0552_ _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_39_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3181_ spi_data_crossing\[31\].A clknet_leaf_7_clock spi_data_crossing\[31\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2305__A2 _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2132_ _0511_ _0108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2063_ _0466_ u1.ordering_complete\[4\] _0462_ _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_35_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3043__CLK clknet_leaf_3_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2965_ _0107_ clknet_leaf_24_clock u1.ordering_complete\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2896_ _0038_ clknet_leaf_2_clock u1.ccr0\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1916_ _0367_ _0036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1847_ u1.col_limit\[6\] _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1778_ _1394_ _1343_ _1344_ _1345_ _1348_ _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__3193__CLK clknet_leaf_30_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1807__A1 _1405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_22_clock_I clknet_2_2__leaf_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output106_I net106 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2232__B2 u1.ordering_complete\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_21_clock clknet_2_3__leaf_clock clknet_leaf_21_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_36_clock clknet_2_0__leaf_clock clknet_leaf_36_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_48_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3066__CLK clknet_leaf_6_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2426__I _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2471__A1 u1.ordering_complete\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2074__I1 u1.ordering_complete\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2750_ _1410_ _0990_ _0991_ _0982_ _0246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_12_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3257__I clknet_leaf_9_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1701_ u1.timer\[19\] _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2681_ _1191_ _0942_ _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2161__I _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2903__CLK clknet_leaf_36_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1632_ u1.timer\[8\] _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1563_ u1.ccr1\[26\] _1180_ _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3302_ net168 net178 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1494_ _1117_ _1118_ _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3233_ net260 clknet_leaf_17_clock net203 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3164_ net55 net239 spi_data_crossing\[23\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2115_ _0471_ u1.ordering_complete\[22\] _0498_ _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2764__C _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3095_ _0229_ clknet_leaf_26_clock u1.timer\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2046_ u0.write_config_n u0.cmd\[21\] u0.cmd\[20\] _0453_ _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_35_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2462__A1 _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2948_ _0090_ clknet_leaf_12_clock u1.ordering_complete\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1568__A3 _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2879_ _0013_ clknet_leaf_7_clock u0.mem_write_n\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input67_I spi_data[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3089__CLK clknet_leaf_29_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2453__A1 _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2926__CLK clknet_leaf_3_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2692__A1 _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2802_ _1282_ _1014_ _1023_ _0266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2747__A2 _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2733_ u1.timer\[20\] _0978_ _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2664_ _1402_ _0927_ _0931_ _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2595_ _0313_ u1.col_limit\[3\] _0316_ u1.col_limit\[2\] _0315_ _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_1615_ _1230_ _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2759__C _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1546_ _1163_ _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout217 u1.row_sel\[4\] net217 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__2380__B1 _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout228 net229 net228 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3231__CLK clknet_leaf_17_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout239 net240 net239 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_1477_ _1100_ u1.ordering_complete\[14\] _1101_ u1.ordering_complete\[13\] _1102_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3216_ net275 clknet_leaf_17_clock net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3147_ spi_data_crossing\[14\].A clknet_leaf_1_clock spi_data_crossing\[14\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3078_ _0006_ clknet_leaf_9_clock u0.run_state\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2949__CLK clknet_leaf_12_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2029_ u1.ccr1\[25\] _0377_ _0443_ _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_23_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1789__A3 _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2038__I1 _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2738__A2 _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1477__A2 u1.ordering_complete\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2674__A1 _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2851__D u0.cmd\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2029__I1 _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2729__A2 _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3104__CLK clknet_leaf_30_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1764__B _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2380_ _0703_ _0682_ _0691_ _0706_ _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_42_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3001_ _0143_ clknet_leaf_17_clock u1.row_col_select\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3270__I net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2087__S _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput6 la_data_in[11] net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__2665__A1 _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2716_ _1303_ _0966_ _0969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2647_ _1216_ _0914_ _1219_ _1202_ _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2578_ _0299_ _0858_ _0859_ spi_data_crossing\[26\].data_sync _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1529_ u0.run_state\[4\] _1151_ _1152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_19_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2656__A1 u1.ccr1\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2408__A1 _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3127__CLK clknet_leaf_36_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output98_I net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2846__D u0.cmd\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2434__I _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1880_ _0330_ _0338_ _0339_ _0028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_30_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2501_ _0796_ _0811_ _0805_ _0810_ _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_2432_ _0752_ _0167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2363_ u1.ordering_timer\[13\] u1.ordering_timer\[12\] _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2294_ _0613_ _0629_ _0631_ _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2638__B2 _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1861__A2 u1.col_limit\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2344__I u1.ordering_timer\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2574__B1 _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput151 net151 io_driver_io_oeb[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput140 net140 io_driver_io_oeb[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput173 net173 mem_address_right[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput162 net162 mem_address_left[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput195 net195 row_col_select[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput184 net184 mem_write_n[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1852__A2 u1.col_limit\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2254__I _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2801__A1 _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_17_clock_I clknet_2_3__leaf_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2332__A3 _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1915__I0 u1.ccr0\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2981_ _0123_ clknet_leaf_16_clock u1.col_limit\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1932_ _0378_ _0041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1863_ u1.col_sel\[6\] u1.col_limit\[6\] _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xinput20 la_data_in[8] net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput31 la_oenb[1] net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput64 spi_data[31] net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput53 spi_data[21] net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_1794_ u1.timer\[25\] _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput42 spi_data[11] net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__1508__I u1.ordering_complete\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2415_ u1.ordering_complete\[19\] _0687_ _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_44_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2346_ _1116_ _0665_ _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2277_ _0614_ _0616_ _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1834__A2 u0.cmd\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1598__B2 _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_hold8_I control_trigger vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1522__A1 _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2185__S _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3020__D _0162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2002__A2 _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1761__A1 _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2200_ u0.cmd\[19\] _0487_ _0350_ _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_26_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3180_ net64 net240 spi_data_crossing\[31\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2131_ _0447_ u1.ordering_complete\[28\] _0489_ _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2062_ _0409_ _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2832__CLK clknet_leaf_10_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1816__A2 _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2982__CLK clknet_leaf_16_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2964_ _0106_ clknet_leaf_24_clock u1.ordering_complete\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1915_ u1.ccr0\[20\] _0366_ _0354_ _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2895_ _0037_ clknet_leaf_3_clock u1.ccr0\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1846_ u1.u1.impulse_gen\[0\] _0308_ _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1777_ _1177_ _1394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_2_clock clknet_2_0__leaf_clock clknet_leaf_2_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1504__A1 _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2069__I _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2329_ _0634_ _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input12_I la_data_in[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1807__A2 _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2232__A2 _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2855__CLK clknet_leaf_16_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2854__D net224 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2471__A2 _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2442__I _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2680_ _0937_ _0942_ _0943_ _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1700_ _1299_ _1316_ _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1631_ u1.ccr1\[8\] _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1982__A1 _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3301_ net167 net177 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1562_ u1.timer\[26\] _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3273__I net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1493_ _1111_ _1112_ _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3232_ net266 clknet_leaf_17_clock net202 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1498__B1 _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3163_ spi_data_crossing\[22\].A clknet_leaf_6_clock spi_data_crossing\[22\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input4_I la_data_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2114_ _0500_ _0101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3094_ _0228_ clknet_leaf_26_clock u1.timer\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3010__CLK clknet_leaf_19_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2045_ u0.cmd\[18\] _0349_ _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2462__A2 _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3160__CLK net239 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2947_ _0089_ clknet_leaf_20_clock u1.ordering_complete\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2878_ _0012_ clknet_leaf_7_clock u0.mem_write_n\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1829_ _0300_ _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2878__CLK clknet_leaf_7_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1489__B1 u1.ordering_timer\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2849__D net289 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3033__CLK clknet_leaf_22_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3183__CLK clknet_leaf_28_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2801_ _0411_ _1021_ _1023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2732_ _0937_ _0979_ _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2663_ _1169_ _1172_ _1175_ _0930_ _1185_ _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_2594_ _0322_ _0326_ _0871_ _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__1707__A1 _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1614_ _1227_ _1231_ _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1545_ u1.timer\[25\] _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xfanout218 u0.cmd\[19\] net218 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2380__A1 _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout229 net233 net229 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3215_ net277 clknet_leaf_17_clock net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1476_ u1.ordering_timer\[13\] _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_41_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3146_ net45 net234 spi_data_crossing\[14\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3077_ _0218_ clknet_leaf_4_clock u0.u11.impulse_gen\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2028_ _0431_ _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_35_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_20_clock clknet_2_3__leaf_clock clknet_leaf_20_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_23_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2082__I _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_35_clock clknet_2_0__leaf_clock clknet_leaf_35_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_40_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output166_I net166 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3056__CLK clknet_leaf_5_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2371__A1 _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3000_ _0142_ clknet_leaf_18_clock u1.row_col_select\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput7 la_data_in[12] net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_40_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2417__A2 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3079__CLK clknet_leaf_12_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2715_ _0945_ _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2646_ _1210_ _1218_ _1205_ _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2577_ _0861_ _0203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2353__A1 _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1528_ _1149_ _1150_ _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2916__CLK clknet_leaf_26_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1459_ _1075_ _1081_ _1083_ _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__1459__A3 _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3129_ spi_data_crossing\[5\].A clknet_leaf_0_clock spi_data_crossing\[5\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2805__I _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2540__I _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_13_clock_I clknet_2_1__leaf_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2715__I _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3221__CLK clknet_leaf_17_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2280__B1 _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2500_ u1.ordering_timer\[27\] _0783_ _0768_ _0784_ _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__2450__I _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2431_ u1.ordering_timer\[21\] _0719_ _0733_ _0751_ _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2335__A1 _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2939__CLK clknet_leaf_4_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2362_ _0634_ _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3281__I net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2293_ u1.ordering_complete\[4\] _0630_ _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_42_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2638__A2 _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2574__B2 spi_data_crossing\[24\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2629_ _0901_ _0900_ _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xoutput130 net130 inverter_select[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__2326__A1 _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput152 net152 io_driver_io_oeb[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput141 net141 io_driver_io_oeb[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput163 net163 mem_address_left[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput174 net174 mem_address_right[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput185 net185 mem_write_n[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA_input42_I spi_data[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput196 net196 row_col_select[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_29_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output129_I net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3244__CLK clknet_leaf_8_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2801__A2 _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2317__A1 _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2857__D net221 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1915__I1 _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2332__A4 _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2980_ _0122_ clknet_leaf_14_clock u1.col_limit\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1931_ u1.ccr0\[25\] _0377_ _0359_ _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_14_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1862_ _0315_ _0323_ _0324_ _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput10 la_data_in[15] net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput21 la_data_in[9] net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3276__I net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput54 spi_data[22] net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__2556__A1 _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput32 la_oenb[2] net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_1793_ _1345_ _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput43 spi_data[12] net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput65 spi_data[3] net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__2308__A1 u1.ordering_timer\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2414_ _0735_ _0736_ _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__3117__CLK clknet_leaf_36_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2345_ _0675_ _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2276_ _1136_ _0615_ _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1598__A2 _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2314__A4 _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2538__A1 _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold50_I u1.row_sel\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2538__B2 spi_data_crossing\[11\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1761__A2 _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2130_ _0508_ _0502_ _0510_ _0107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2061_ _0465_ _0083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3211__D _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2077__I0 _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2963_ _0105_ clknet_leaf_20_clock u1.ordering_complete\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1914_ u0.cmd\[4\] _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_33_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2894_ _0036_ clknet_leaf_2_clock u1.ccr0\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1845_ u1.u1.impulse_gen\[1\] _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_11_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1776_ _1330_ _1331_ _1342_ _1386_ _1392_ _1393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__1752__A2 u1.ccr0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2328_ _0661_ _0154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1504__A2 u1.ordering_complete\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2259_ _1403_ _0595_ _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_26_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2465__B1 _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1807__A3 _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3121__D spi_data_crossing\[1\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output196_I net196 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2299__A3 _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2196__S _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1431__A1 _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1630_ u1.timer\[9\] _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1783__B _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3300_ net166 net176 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1561_ _1176_ u1.timer\[27\] _1178_ u1.timer\[26\] _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_45_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1492_ _1116_ u1.ordering_complete\[10\] _1109_ u1.ordering_complete\[9\] _1117_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3231_ net284 clknet_leaf_17_clock net201 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1498__A1 _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3162_ net54 net239 spi_data_crossing\[22\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1498__B2 u1.ordering_complete\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2113_ _0468_ u1.ordering_complete\[21\] _0498_ _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_27_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3093_ _0227_ clknet_leaf_26_clock u1.timer\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2044_ u0.cmd\[16\] _0394_ _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__2119__B _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2946_ _0088_ clknet_leaf_19_clock u1.ordering_complete\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2877_ _0011_ clknet_leaf_12_clock u0.timer_enable vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1828_ _0296_ _0301_ _0013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1759_ _1363_ u1.ccr0\[1\] _1366_ _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1489__A1 u1.ordering_timer\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1489__B2 _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1712__I u1.ccr0\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output209_I net209 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1661__A1 _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2213__I0 _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2972__CLK clknet_leaf_9_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2718__I _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_2_1__f_clock clknet_0_clock clknet_2_1__leaf_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_1_clock clknet_2_0__leaf_clock clknet_leaf_1_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_32_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2800_ _1286_ _1014_ _1022_ _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2731_ _1224_ _0978_ _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_8_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2662_ u1.ccr1\[28\] _1173_ u1.ccr1\[27\] _1349_ _1179_ _0929_ _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__2204__I0 _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3284__I net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2593_ _0312_ _0324_ _0870_ _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1613_ u1.ccr1\[23\] _1228_ u1.ccr1\[22\] _1229_ u1.ccr1\[21\] _1230_ _1231_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_1544_ _1043_ _1162_ _0007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1707__A2 _1320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2380__A2 _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout219 u0.cmd\[15\] net219 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3214_ net267 clknet_leaf_17_clock net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1475_ u1.ordering_timer\[14\] _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_45_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2628__I net216 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3145_ spi_data_crossing\[13\].A clknet_leaf_1_clock spi_data_crossing\[13\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3076_ _0217_ clknet_leaf_5_clock u0.u11.impulse_gen\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2027_ _0442_ _0072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2845__CLK clknet_leaf_15_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2929_ _0071_ clknet_leaf_2_clock u1.ccr1\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input72_I spi_data_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2995__CLK clknet_leaf_16_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2371__A2 _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output159_I net159 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1442__I u1.ordering_complete\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2273__I _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3000__CLK clknet_leaf_18_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput8 la_data_in[13] net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__1873__A1 _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3279__I net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2868__CLK clknet_leaf_11_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1625__A1 u1.ccr1\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2714_ _0958_ _0966_ _0967_ _0234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2645_ _0912_ _1198_ _1201_ _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_12_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2576_ u0.cmd\[25\] _0858_ _0859_ spi_data_crossing\[25\].data_sync _0861_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1527_ u0.run_state\[5\] _1044_ u0.run_state\[1\] _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_45_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1458_ u1.ordering_timer\[31\] _1073_ _1082_ _1078_ _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_19_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3128_ net67 net227 spi_data_crossing\[5\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3059_ _0201_ clknet_leaf_6_clock u0.cmd\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1616__A1 u1.ccr1\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3023__CLK clknet_leaf_21_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3173__CLK clknet_leaf_7_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2280__A1 u1.ordering_timer\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2430_ u1.ordering_complete\[21\] _0750_ _0609_ _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_29_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2361_ _0690_ _0158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2379__S _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2292_ _0608_ _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2178__I _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_34_clock clknet_2_0__leaf_clock clknet_leaf_34_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_17_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3046__CLK clknet_leaf_1_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3196__CLK clknet_leaf_24_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2574__A2 _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1782__B1 _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput120 net120 data_out_right[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_2628_ net216 _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput131 net131 inverter_select[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput142 net142 io_driver_io_oeb[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput164 net164 mem_address_left[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput175 net175 mem_address_right[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput186 net186 mem_write_n[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_2559_ _0850_ _0196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput153 net153 io_driver_io_oeb[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput197 net197 row_col_select[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_47_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input35_I la_oenb[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2262__A1 _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2551__I _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3069__CLK clknet_leaf_9_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1930_ u0.cmd\[9\] _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2253__A1 _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1861_ _0311_ u1.col_limit\[5\] _0314_ u1.col_limit\[4\] _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_14_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout222_I u0.cmd\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput11 la_data_in[16] net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput22 la_oenb[0] net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__2906__CLK clknet_leaf_30_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput55 spi_data[23] net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_7_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput33 la_oenb[3] net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_1792_ _1406_ _1407_ _1408_ _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xinput44 spi_data[13] net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_6_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput66 spi_data[4] net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2413_ _1064_ _0728_ _0724_ _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_2344_ u1.ordering_timer\[11\] _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2275_ _1138_ _0599_ _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3119__D spi_data_crossing\[0\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3211__CLK clknet_leaf_33_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2483__A1 _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2235__A1 _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2929__CLK clknet_leaf_2_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2710__A2 _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2060_ _0464_ u1.ordering_complete\[3\] _0462_ _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_35_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2077__I1 _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2962_ _0104_ clknet_leaf_20_clock u1.ordering_complete\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1913_ _1319_ _0360_ _0365_ _0035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2893_ _0035_ clknet_leaf_2_clock u1.ccr0\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1844_ _0307_ net33 _0024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1775_ _1337_ _1391_ _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3234__CLK clknet_leaf_7_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2327_ _0654_ _0655_ _0635_ _0660_ _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2258_ u1.ordering_timer\[1\] _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2189_ _0546_ _0130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2465__A1 _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3107__CLK clknet_leaf_31_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1431__A2 u1.ordering_complete\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1560_ u1.ccr1\[26\] _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1491_ u1.ordering_timer\[10\] _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1990__I0 u1.ccr1\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3230_ net264 clknet_leaf_17_clock net200 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1498__A2 u1.ordering_complete\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3161_ spi_data_crossing\[21\].A clknet_leaf_6_clock spi_data_crossing\[21\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2695__A1 _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2112_ _0499_ _0100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3092_ _0226_ clknet_leaf_25_clock u1.timer\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2043_ _0451_ _0079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2945_ _0087_ clknet_leaf_19_clock u1.ordering_complete\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2876_ _0022_ clknet_leaf_6_clock u0.write_config_n vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1827_ _0299_ _1149_ _0300_ _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_11_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1758_ _1299_ _1316_ _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1689_ _1303_ _1304_ _1305_ _1254_ _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1489__A2 _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2686__A1 _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2438__A1 _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output104_I net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1661__A2 _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2374__B1 _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2677__A1 _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1652__A2 _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2730_ _0968_ _0977_ _0978_ _0239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_8_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2661_ _0928_ _1181_ _1183_ _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1612_ u1.timer\[21\] _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2592_ net226 _0321_ _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1543_ u0.run_state\[3\] _1144_ _1161_ _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1474_ _1096_ _1097_ u1.ordering_timer\[14\] _1098_ _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3213_ _0000_ clknet_leaf_32_clock control_trigger vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3144_ net44 net231 spi_data_crossing\[13\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3075_ _0216_ clknet_leaf_11_clock u1.row_sel\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2026_ u1.ccr1\[24\] _0375_ _0432_ _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_17_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2928_ _0070_ clknet_leaf_31_clock u1.ccr1\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2859_ net219 clknet_leaf_16_clock net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input65_I spi_data[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2659__A1 _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2131__I0 _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2198__I0 _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput9 la_data_in[14] net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__1873__A2 _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2122__I0 _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1625__A2 _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2822__A1 net220 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2713_ _1300_ _0963_ _1254_ _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_10_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2644_ _1200_ _1188_ _1196_ _1190_ _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2575_ _0860_ _0202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1526_ u0.cmd\[27\] _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_45_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1457_ u1.ordering_timer\[30\] _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3127_ spi_data_crossing\[4\].A clknet_leaf_36_clock spi_data_crossing\[4\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3058_ _0200_ clknet_leaf_6_clock u0.cmd\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2113__I0 _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1616__A2 _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2813__A1 net224 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2009_ _0427_ _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_24_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2962__CLK clknet_leaf_20_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1552__A1 u1.ccr1\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_0_clock clknet_2_0__leaf_clock clknet_leaf_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__2549__I _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2280__A2 _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2032__A2 _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1791__A1 _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2360_ u1.ordering_timer\[12\] _0682_ _0662_ _0689_ _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_29_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2291_ _1122_ _0628_ _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_49_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2835__CLK clknet_leaf_10_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2985__CLK clknet_leaf_16_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2023__A2 _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput110 net110 data_out_left[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__1782__A1 _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput121 net121 data_out_right[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_2627_ _0890_ _0899_ _0900_ _0214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
Xoutput132 net132 inverter_select[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput143 net143 io_driver_io_oeb[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput165 net165 mem_address_left[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput176 net176 mem_address_right[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_2558_ u0.cmd\[18\] _0845_ _0847_ spi_data_crossing\[18\].data_sync _0850_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput154 net154 io_driver_io_oeb[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput187 net187 mem_write_n[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput198 net198 row_col_select[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_1509_ u1.ordering_complete\[1\] _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2489_ _0800_ _0801_ _0714_ _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input28_I la_oenb[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2247__C1 _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2262__A2 _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1448__I u1.ordering_complete\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output96_I net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2858__CLK clknet_leaf_16_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1525__A1 _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1828__A2 _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1911__I u0.cmd\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1860_ _0313_ u1.col_limit\[3\] _0316_ u1.col_limit\[2\] _0320_ _0322_ _0323_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
Xinput12 la_data_in[17] net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_1791_ _1272_ _1295_ _1248_ _1250_ _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_35_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput34 la_oenb[4] net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput23 la_oenb[10] net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput45 spi_data[14] net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput56 spi_data[24] net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput67 spi_data[5] net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__1764__A1 _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1516__A1 _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2412_ u1.ordering_timer\[18\] _0723_ _0583_ _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2343_ _0674_ _0156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_42_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2274_ _1138_ _0599_ u1.ordering_timer\[2\] _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_42_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3013__CLK clknet_leaf_19_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2492__A2 _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3163__CLK clknet_leaf_6_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1989_ _1247_ _0414_ _0419_ _0057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2099__I _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2827__I _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2483__A2 _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2562__I _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_33_clock clknet_2_0__leaf_clock clknet_leaf_33_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__1906__I _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3036__CLK clknet_leaf_3_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2737__I _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3186__CLK clknet_leaf_33_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2961_ _0103_ clknet_leaf_21_clock u1.ordering_complete\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1912_ _0364_ _0362_ _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1985__A1 u0.cmd\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2892_ _0034_ clknet_leaf_2_clock u1.ccr0\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1843_ net15 _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1737__A1 _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1774_ _1333_ _1390_ _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1737__B2 u1.timer\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2326_ _0643_ _0657_ _0659_ _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2257_ _0565_ _0598_ _0146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_38_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2188_ _0466_ u1.inverter_select\[4\] _0545_ _0546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_26_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2465__A2 _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2382__I _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3059__CLK clknet_leaf_6_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1726__I u1.ccr0\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1461__I u1.ordering_complete\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1719__A1 _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2392__A1 _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1490_ _1109_ _1110_ _1111_ _1112_ _1114_ _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_4_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1990__I1 _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3160_ net53 net239 spi_data_crossing\[21\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2111_ _0466_ u1.ordering_complete\[20\] _0498_ _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3091_ _0225_ clknet_leaf_25_clock u1.timer\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold1 latch_data net243 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XANTENNA__2467__I u1.ordering_timer\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2042_ u1.ccr1\[31\] _0390_ _0431_ _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_47_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2447__A2 _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1655__B1 u1.ccr1\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3298__I net164 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2944_ _0086_ clknet_leaf_19_clock u1.ordering_complete\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2875_ u0.latch_cmd clknet_leaf_4_clock u0.update_cmd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1826_ u0.cmd\[31\] _0297_ _0300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3201__CLK clknet_leaf_23_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1757_ _1317_ _1342_ _1373_ _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1688_ u1.ccr0\[14\] _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2919__CLK clknet_leaf_27_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2135__A1 u0.cmd\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2309_ u1.ordering_complete\[6\] _0630_ _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2686__A2 _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3289_ net155 net154 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input10_I la_data_in[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2374__A1 _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2429__A2 _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1637__B1 _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3224__CLK clknet_leaf_16_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2660_ u1.ccr1\[25\] _1164_ u1.ccr1\[24\] _1166_ _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1611_ u1.timer\[22\] _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2591_ _0869_ _0209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1542_ _1159_ _1045_ _1150_ _1160_ _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_5_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1473_ u1.ordering_complete\[14\] _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_45_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3212_ _0002_ clknet_leaf_34_clock latch_data vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input2_I io_latch_data_in vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2668__A2 _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3143_ spi_data_crossing\[12\].A clknet_leaf_0_clock spi_data_crossing\[12\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3074_ _0215_ clknet_leaf_10_clock u1.row_sel\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2025_ _1225_ _0435_ _0441_ _0071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2927_ _0069_ clknet_leaf_2_clock u1.ccr1\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2858_ net220 clknet_leaf_16_clock net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1809_ net16 net3 net34 _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2789_ _0392_ _1015_ _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input58_I spi_data[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2108__A1 _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2891__CLK clknet_leaf_2_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3143__D spi_data_crossing\[12\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3247__CLK clknet_leaf_8_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2131__I1 u1.ordering_complete\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1914__I u0.cmd\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2011__S _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2822__A2 _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2586__B2 spi_data_crossing\[29\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2586__A1 u0.cmd\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2712_ _1254_ _1300_ _1262_ _0961_ _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_2643_ u1.ccr1\[7\] _1193_ _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2574_ u0.cmd\[24\] _0858_ _0859_ spi_data_crossing\[24\].data_sync _0860_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1525_ _1043_ _1148_ _0009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_45_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1456_ _1077_ _1080_ _1081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3126_ net66 net227 spi_data_crossing\[4\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3057_ _0199_ clknet_leaf_5_clock u0.cmd\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__2113__I1 u1.ordering_complete\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2008_ _0430_ _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2390__I _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output164_I net164 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2501__A1 _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2804__A2 _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2568__A1 u0.cmd\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1918__I1 _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1543__A2 _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2740__A1 _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2290_ u1.ordering_timer\[0\] u1.ordering_timer\[1\] u1.ordering_timer\[3\] u1.ordering_timer\[2\]
+ _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_1_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1819__I u0.cmd\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput100 net100 data_out_left[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_2626_ net217 _0897_ _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1782__A2 u1.ccr0\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput122 net122 data_out_right[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput111 net111 data_out_right[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput133 net133 inverter_select[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_12_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput177 net177 mem_address_right[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput166 net166 mem_address_left[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_47_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2557_ _0849_ _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput155 net155 io_driver_io_oeb[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput144 net144 io_driver_io_oeb[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__2731__A1 _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3092__CLK clknet_leaf_25_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput199 net199 row_col_select[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput188 net188 mem_write_n[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_1508_ u1.ordering_complete\[0\] _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2488_ _1076_ _0796_ _1093_ _0790_ _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_1439_ u1.ordering_timer\[19\] _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_46_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1837__A3 _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3109_ _0243_ clknet_leaf_31_clock u1.timer\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2247__B1 u1.ordering_timer\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2247__C2 _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1470__A1 _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2089__I0 _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2789__A1 _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput13 la_data_in[1] net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_11_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1790_ _1206_ _1208_ _1214_ _1203_ _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
Xinput46 spi_data[15] net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput35 la_oenb[5] net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput24 la_oenb[11] net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput57 spi_data[25] net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput68 spi_data[6] net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_13_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2411_ _0608_ _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2342_ u1.ordering_timer\[10\] _0655_ _0662_ _0673_ _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2273_ _0612_ _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2952__CLK clknet_leaf_3_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1549__I u1.timer\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1452__A1 _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1452__B2 u1.ordering_complete\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1988_ u0.cmd\[9\] _0418_ _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2609_ u1.row_sel\[6\] _0526_ _0524_ net216 _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2704__A1 _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input40_I spi_data[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1994__A2 _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2794__I1 _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2975__CLK clknet_leaf_11_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1682__A1 _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2960_ _0102_ clknet_leaf_20_clock u1.ordering_complete\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1809__I0 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1911_ u0.cmd\[3\] _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2891_ _0033_ clknet_leaf_2_clock u1.ccr0\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1842_ _0306_ _0004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1773_ _1338_ _1389_ _1335_ _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_48_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3236__D u0.cmd\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2325_ _1112_ _0658_ _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2256_ _1139_ _0597_ _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_38_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2187_ _0539_ _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2848__CLK clknet_leaf_16_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2998__CLK clknet_leaf_18_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2573__I _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3003__CLK clknet_leaf_18_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1917__I u0.cmd\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3153__CLK clknet_leaf_5_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold2 u0.mem_write_n\[9\] net244 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_2110_ _0491_ _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3090_ _0224_ clknet_leaf_23_clock u1.timer\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2041_ _0450_ _0078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1655__B2 _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2943_ _0085_ clknet_leaf_14_clock u1.ordering_complete\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2874_ _0031_ clknet_leaf_16_clock u1.col_sel\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1825_ u0.cmd\[26\] _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1756_ _1362_ _1372_ _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1687_ u1.ccr0\[15\] _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_48_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2135__A2 _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2308_ u1.ordering_timer\[6\] _0636_ _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3288_ net153 net152 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2239_ _1210_ _0580_ _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_32_clock clknet_2_0__leaf_clock clknet_leaf_32_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_14_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3026__CLK clknet_leaf_20_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3176__CLK net238 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2374__A2 _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1472__I u1.ordering_complete\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2126__A2 _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1885__A1 _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2677__A3 _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1637__B2 _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1610_ u1.timer\[23\] _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2590_ _1040_ _0864_ _0865_ spi_data_crossing\[31\].data_sync _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1541_ u0.cmd\[27\] _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1472_ u1.ordering_complete\[15\] _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3211_ _0003_ clknet_leaf_33_clock reset_n vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3142_ net43 net231 spi_data_crossing\[12\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1876__A1 _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3073_ _0214_ clknet_leaf_10_clock u1.row_sel\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1628__A1 _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2024_ _0373_ _0436_ _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3049__CLK clknet_leaf_4_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2053__A1 _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3199__CLK clknet_leaf_31_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2926_ _0068_ clknet_leaf_3_clock u1.ccr1\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2857_ net221 clknet_leaf_15_clock net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1808_ _1401_ _1403_ _0289_ _0023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__2356__A2 _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2788_ _1012_ _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1739_ _1348_ _1350_ _1354_ _1355_ _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__2108__A2 _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1867__A1 _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output207_I net207 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2044__A1 u0.cmd\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2595__A2 u1.col_limit\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1930__I u0.cmd\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2283__A1 u1.ordering_complete\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout238_I net239 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2909__CLK clknet_leaf_22_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2711_ _0935_ _0965_ _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_13_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2642_ _1255_ _0909_ _1260_ _1264_ _0910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2573_ _0846_ _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2202__S _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1524_ u0.cmd\[28\] u0.run_state\[2\] _1147_ u0.run_state\[5\] _1148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_5_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1455_ u1.ordering_timer\[30\] _1078_ u1.ordering_timer\[29\] _1079_ _1080_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_28_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3125_ spi_data_crossing\[3\].A clknet_leaf_36_clock spi_data_crossing\[3\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3056_ _0198_ clknet_leaf_5_clock u0.cmd\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_2007_ u1.ccr1\[17\] _0400_ _0428_ _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2671__I _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2909_ _0051_ clknet_leaf_22_clock u1.ccr1\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input70_I spi_data[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2620__B u1.row_sel\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3214__CLK clknet_leaf_17_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2501__A2 _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1750__I _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1776__B1 _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1791__A3 _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2040__I1 _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2881__CLK clknet_leaf_8_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3239__D u0.cmd\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2625_ net217 _0897_ _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xoutput101 net101 data_out_left[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_12_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput112 net112 data_out_right[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput123 net123 data_out_right[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__3237__CLK clknet_leaf_7_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput134 net134 inverter_select[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput167 net167 mem_address_left[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_2556_ _0348_ _0845_ _0847_ spi_data_crossing\[17\].data_sync _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput156 net156 io_driver_io_oeb[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput145 net145 io_driver_io_oeb[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput178 net178 mem_address_right[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput189 net189 mem_write_n[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_1507_ _1127_ _1130_ _1131_ _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_2487_ u1.ordering_timer\[28\] _0791_ u1.ordering_timer\[29\] _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_25_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1438_ u1.ordering_timer\[19\] _1058_ _1059_ _1060_ _1062_ _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XANTENNA__2666__I _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2495__A1 _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3108_ _0242_ clknet_leaf_31_clock u1.timer\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3039_ _0181_ clknet_leaf_4_clock u0.cmd\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2247__A1 u1.ordering_timer\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1470__A2 _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2722__A2 _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2486__A1 _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2089__I1 u1.ordering_complete\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2253__A4 _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput14 la_data_in[2] net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput36 la_oenb[6] net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput25 la_oenb[12] net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput58 spi_data[26] net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput47 spi_data[16] net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput69 spi_data[7] net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_48_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2410_ _0634_ _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2341_ _0670_ _0671_ _0672_ _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2713__A2 _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2272_ _0607_ _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1452__A2 u1.ordering_complete\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1987_ _0397_ _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2401__A1 _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2608_ _0524_ net216 _0521_ net217 _0885_ _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_2539_ _0837_ _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input33_I la_oenb[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2468__A1 _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1475__I u1.ordering_timer\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2459__A1 _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1682__A2 u1.ccr0\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3082__CLK clknet_leaf_4_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1809__I1 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2631__A1 net216 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1910_ _1320_ _0360_ _0363_ _0034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2890_ _0032_ clknet_leaf_3_clock u1.ccr0\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1841_ _0304_ u0.run_state\[2\] _1155_ _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_8_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout220_I u0.cmd\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1772_ _1323_ _1325_ _1387_ _1388_ _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2698__A1 _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2324_ _0596_ _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2255_ _0596_ _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2186_ _0544_ _0129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2120__S _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2689__A1 u1.timer\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2942__CLK clknet_leaf_14_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1933__I _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold3 u0.mem_write_n\[7\] net245 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_48_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2040_ u1.ccr1\[30\] _0388_ _0443_ _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_35_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1655__A2 _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2942_ _0084_ clknet_leaf_14_clock u1.ordering_complete\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2604__A1 u1.row_limit\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2604__B2 _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2873_ _0030_ clknet_leaf_16_clock u1.col_sel\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2713__B _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1824_ _0296_ _0298_ _0012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2368__B1 _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1755_ _1366_ _1368_ _1371_ _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__2004__I _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1686_ u1.timer\[15\] _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2307_ _0612_ _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3287_ net151 net150 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1894__A2 u0.cmd\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2238_ _1205_ _1216_ _1217_ _1220_ _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__2143__I0 _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2169_ _0464_ u1.col_limit\[3\] _0529_ _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1646__A2 u1.timer\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2965__CLK clknet_leaf_24_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2115__S _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output187_I net187 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1637__A2 u1.timer\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3120__CLK net229 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1540_ u0.run_state\[6\] _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_8_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1471_ u1.ordering_timer\[15\] _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1663__I _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2838__CLK clknet_leaf_15_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3210_ _0279_ clknet_leaf_35_clock net137 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3141_ spi_data_crossing\[11\].A clknet_leaf_0_clock spi_data_crossing\[11\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1876__A2 _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3072_ _0213_ clknet_leaf_10_clock u1.row_sel\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2988__CLK clknet_leaf_18_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2023_ _1226_ _0435_ _0440_ _0070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2053__A2 _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2925_ _0067_ clknet_leaf_30_clock u1.ccr1\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2856_ net222 clknet_leaf_16_clock net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1807_ _1405_ _1409_ _0280_ _0288_ _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_15_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2787_ _1013_ _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1738_ _1171_ u1.ccr0\[31\] u1.ccr0\[24\] _1166_ _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_46_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1669_ u1.ccr0\[4\] _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_24_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2816__A1 net223 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output102_I net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_7_clock_I clknet_2_1__leaf_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3143__CLK clknet_leaf_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2807__A1 _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2283__A2 _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2710_ _1258_ _0963_ _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_12_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2641_ _1252_ _1303_ _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2572_ _0844_ _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_31_clock clknet_2_0__leaf_clock clknet_leaf_31_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1523_ control_trigger_sync\[0\] control_trigger control_trigger_sync\[1\] _1147_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1454_ u1.ordering_complete\[29\] _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_45_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1849__A2 u1.col_limit\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3016__CLK clknet_leaf_14_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3124_ net65 net227 spi_data_crossing\[3\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3055_ _0197_ clknet_leaf_5_clock u0.cmd\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2006_ _0429_ _0064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2908_ _0050_ clknet_leaf_22_clock u1.ccr1\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2839_ net295 clknet_leaf_10_clock net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input63_I spi_data[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1517__B _1140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2399__I _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2017__A2 _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1776__B2 _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1791__A4 _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3039__CLK clknet_leaf_4_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3189__CLK clknet_leaf_35_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1700__A1 _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2256__A2 _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2624_ _0890_ _0897_ _0898_ _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__2213__S _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput113 net113 data_out_right[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput124 net124 data_out_right[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput102 net102 data_out_left[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput168 net168 mem_address_left[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput135 net135 inverter_select[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_2555_ _0848_ _0194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput157 net157 io_driver_io_oeb[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput146 net146 io_driver_io_oeb[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput179 net179 mem_address_right[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_1506_ _1125_ u1.ordering_complete\[6\] _1121_ u1.ordering_complete\[5\] _1131_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_2486_ _0796_ _0710_ _0799_ _0174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1437_ u1.ordering_timer\[17\] _1061_ u1.ordering_timer\[16\] _1060_ _1062_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_29_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2495__A2 _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3107_ _0241_ clknet_leaf_31_clock u1.timer\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3038_ _0180_ clknet_leaf_3_clock u0.cmd\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1470__A3 _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1758__A1 _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2486__A2 _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1997__A1 net221 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput15 la_data_in[3] net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput37 la_oenb[7] net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput26 la_oenb[13] net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput59 spi_data[27] net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput48 spi_data[17] net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_7_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2340_ u1.ordering_complete\[10\] _0658_ _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_46_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2271_ _0611_ _0147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_2_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2767__I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2208__S _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_34_clock_I clknet_2_0__leaf_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1988__A1 u0.cmd\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3204__CLK clknet_leaf_23_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1986_ _1249_ _0414_ _0417_ _0056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_18_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2401__A2 _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2607_ u1.row_limit\[4\] _0876_ u1.row_limit\[3\] _0877_ _0884_ _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__2165__A1 _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2538_ _0382_ _0832_ _0833_ spi_data_crossing\[11\].data_sync _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1581__I u1.ccr1\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1912__A1 _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2469_ _0768_ _0784_ _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_29_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input26_I la_oenb[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3301__I net167 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1979__A1 _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1491__I u1.ordering_timer\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2871__CLK clknet_leaf_15_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2459__A2 _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1667__B1 _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3227__CLK clknet_leaf_17_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1840_ _0304_ _1153_ _0301_ _0021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_37_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1771_ _1336_ _1334_ _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2323_ _1111_ _0656_ _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2254_ _0595_ _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2185_ _0464_ u1.inverter_select\[3\] _0540_ _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_38_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2622__A2 _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2386__A1 _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1576__I u1.timer\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1969_ _1215_ _0403_ _0406_ _0050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2138__A1 _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2689__A2 u1.timer\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2894__CLK clknet_leaf_2_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2310__A1 _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2377__A1 _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2129__A1 u0.cmd\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2110__I _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold4 u0.mem_write_n\[8\] net246 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_0_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2301__A1 _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2941_ _0083_ clknet_leaf_14_clock u1.ordering_complete\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2872_ _0029_ clknet_leaf_14_clock u1.col_sel\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1823_ u0.cmd\[31\] u0.cmd\[26\] u0.cmd\[27\] _0297_ _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__2368__A1 u1.ordering_timer\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1754_ _1364_ u1.ccr0\[0\] _1369_ _1370_ _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__2221__S _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1685_ _1300_ _1301_ _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_48_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2306_ _0642_ _0151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_38_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3286_ net149 net138 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1894__A3 u0.cmd\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2237_ _1187_ _1235_ _1245_ _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_22_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2168_ _0319_ _0530_ _0534_ _0121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2099_ _0488_ _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2359__A1 _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2131__S _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_3_clock_I clknet_2_1__leaf_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3072__CLK clknet_leaf_10_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3173__D spi_data_crossing\[27\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2295__B1 _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2105__I _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2770__A1 _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1470_ _1084_ _1090_ _1092_ _1094_ _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_45_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2522__A1 _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2522__B2 spi_data_crossing\[4\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3140_ net42 net230 spi_data_crossing\[11\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3071_ _0212_ clknet_leaf_9_clock u1.row_sel\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2022_ _0370_ _0436_ _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2924_ _0066_ clknet_leaf_3_clock u1.ccr1\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2855_ net223 clknet_leaf_16_clock net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1806_ _0284_ _0287_ _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2015__I _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2786_ _1012_ _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2761__A1 u1.timer\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3095__CLK clknet_leaf_26_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1737_ _1351_ _1352_ _1353_ u1.timer\[30\] _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1668_ _1193_ u1.ccr0\[7\] u1.ccr0\[4\] _1194_ _1284_ _1285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_1599_ _1207_ u1.ccr1\[0\] _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3269_ net88 net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2932__CLK clknet_2_0__leaf_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2796__S _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2036__S _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2640_ _1274_ _1251_ _1275_ _0907_ _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_16_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2571_ _0857_ _0201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1522_ _1043_ _1146_ _0010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2743__A1 _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1453_ u1.ordering_complete\[30\] _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2955__CLK clknet_leaf_3_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3123_ spi_data_crossing\[2\].A clknet_leaf_36_clock spi_data_crossing\[2\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3054_ _0196_ clknet_leaf_5_clock u0.cmd\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2005_ u1.ccr1\[16\] _0392_ _0428_ _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_24_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2274__A3 u1.ordering_timer\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1482__A1 _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2431__B1 _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2907_ _0049_ clknet_leaf_30_clock u1.ccr1\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2838_ net268 clknet_leaf_15_clock net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2769_ net10 _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2734__A1 u1.timer\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input56_I spi_data[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_29_clock_I clknet_2_2__leaf_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3304__I net170 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3110__CLK clknet_leaf_33_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2422__B1 _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2978__CLK clknet_leaf_11_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1528__A2 _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2725__A1 _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1464__A1 _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2623_ u1.row_sel\[3\] _0895_ _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_12_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput103 net103 data_out_left[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput114 net114 data_out_right[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput125 net125 data_out_right[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__1519__A2 _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2554_ _0393_ _0845_ _0847_ spi_data_crossing\[16\].data_sync _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2716__A1 _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput136 net136 inverter_select[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_1505_ _1128_ u1.ordering_complete\[3\] _1122_ u1.ordering_complete\[4\] _1129_ _1130_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
Xoutput158 net158 io_latch_data_oeb vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput147 net147 io_driver_io_oeb[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput169 net169 mem_address_left[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_2485_ u1.ordering_complete\[28\] _0720_ _0604_ _0798_ _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA_clkbuf_leaf_30_clock_I clknet_2_0__leaf_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1436_ u1.ordering_complete\[17\] _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__3133__CLK clknet_leaf_5_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3106_ _0240_ clknet_leaf_31_clock u1.timer\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3037_ _0179_ clknet_leaf_3_clock u0.cmd\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1455__A1 u1.ordering_timer\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2007__I0 u1.ccr1\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2707__A1 _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output162_I net162 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_30_clock clknet_2_0__leaf_clock clknet_leaf_30_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__1997__A2 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3006__CLK clknet_leaf_12_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput16 la_data_in[4] net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput27 la_oenb[14] net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_11_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput49 spi_data[18] net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput38 la_oenb[8] net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_13_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1952__I u0.cmd\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2270_ _0599_ _0602_ _0605_ _0610_ _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_42_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2783__I u1.ccr0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1437__B2 _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1988__A2 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1985_ u0.cmd\[8\] _0412_ _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2606_ _0880_ _0882_ _0883_ _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2165__A2 _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2537_ _0836_ _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2468_ _0773_ _0760_ u1.ordering_timer\[22\] _0748_ _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__1912__A2 _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1419_ control_trigger_sync\[0\] control_trigger control_trigger_sync\[1\] _1044_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_29_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2399_ _0723_ _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2468__A3 u1.ordering_timer\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input19_I la_data_in[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1428__B2 u1.ordering_complete\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1979__A2 _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3029__CLK clknet_leaf_24_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3179__CLK clknet_leaf_6_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1600__A1 u1.ccr1\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1667__B2 _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2092__A1 _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2219__I0 _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1770_ _1323_ _1326_ _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2322_ _0648_ _0649_ _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2253_ _1212_ _0578_ _0582_ _0594_ _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_2184_ _0543_ _0128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1658__A1 u1.ccr1\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2219__S _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2083__A1 net224 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1830__A1 u0.cmd\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2386__A2 _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1968_ _0404_ _0405_ _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1899_ u1.ccr0\[16\] _0346_ _0354_ _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_1_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2138__A2 _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2689__A3 _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3312__I net209 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1821__A1 u0.cmd\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2377__A2 _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2598__I net217 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2129__A2 _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1888__A1 _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold27_I u0.cmd\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold5 u0.mem_write_n\[4\] net247 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_0_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2940_ _0082_ clknet_leaf_13_clock u1.ordering_complete\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2871_ _0028_ clknet_leaf_15_clock u1.col_sel\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1822_ _0295_ u0.update_cmd _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2368__A2 _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1753_ _1204_ u1.ccr0\[2\] _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2502__S _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1684_ u1.ccr0\[13\] _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1879__A1 u1.col_sel\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3285_ net101 net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2305_ u1.ordering_timer\[5\] _0627_ _0635_ _0641_ _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1894__A4 u0.cmd\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2236_ _0566_ _0577_ _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_26_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2167_ _0404_ _0531_ _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2098_ _0489_ _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2861__CLK clknet_leaf_5_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3307__I net204 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3217__CLK clknet_leaf_16_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3070_ _0211_ clknet_leaf_9_clock u1.row_sel\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2021_ _0439_ _0069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2791__I _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2884__CLK clknet_leaf_8_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2923_ _0065_ clknet_leaf_2_clock u1.ccr1\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2854_ net224 clknet_leaf_16_clock net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1805_ _0285_ _0286_ u1.timer\[21\] u1.timer\[20\] _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_2785_ _1011_ _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1736_ u1.ccr0\[30\] _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_49_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1667_ _1280_ _1281_ _1282_ _1283_ _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1598_ _1213_ _1214_ _1215_ _1203_ _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_24_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3268_ net87 net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2219_ _0476_ u1.row_col_select\[8\] _0552_ _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_27_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3199_ _0269_ clknet_leaf_31_clock u1.ccr0\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_25_clock_I clknet_2_2__leaf_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output192_I net192 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2650__B _0910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3184__D _0254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2570_ u0.cmd\[23\] _0852_ _0853_ spi_data_crossing\[23\].data_sync _0857_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1521_ u0.run_state\[6\] _1045_ _1145_ u0.run_state\[3\] _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_5_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1452_ _1076_ u1.ordering_complete\[29\] _1071_ u1.ordering_complete\[28\] _1077_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__2786__I _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3122_ net62 net229 spi_data_crossing\[2\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3053_ _0195_ clknet_leaf_5_clock u0.cmd\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2259__A1 _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2004_ _0427_ _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1482__A2 u1.ordering_complete\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3062__CLK clknet_leaf_8_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2431__A1 u1.ordering_timer\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2906_ _0048_ clknet_leaf_30_clock u1.ccr1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2837_ net276 clknet_leaf_10_clock net209 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2768_ _1002_ net29 _0253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2699_ _0946_ _0956_ _0957_ _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1719_ _1236_ u1.ccr0\[17\] _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input49_I spi_data[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2498__A1 _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output205_I net205 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2670__A1 _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3179__D spi_data_crossing\[30\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3085__CLK clknet_leaf_35_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1464__A2 u1.ordering_complete\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2413__A1 _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout236_I net241 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2622_ u1.row_sel\[3\] _0895_ _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2922__CLK clknet_leaf_2_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput115 net115 data_out_right[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput104 net104 data_out_left[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_2553_ _0846_ _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1519__A3 _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2716__A2 _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput126 net126 data_out_right[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_1504_ _1124_ u1.ordering_complete\[7\] _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xoutput159 net159 io_reset_n_oeb vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput137 net137 io_control_trigger_oeb vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput148 net148 io_driver_io_oeb[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_2484_ _0597_ _0797_ _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1435_ u1.ordering_complete\[16\] _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_29_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3105_ _0239_ clknet_leaf_31_clock u1.timer\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3036_ _0178_ clknet_leaf_3_clock u0.cmd\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1455__A2 _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2007__I1 _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2707__A2 _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2643__A1 u1.ccr1\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2945__CLK clknet_leaf_19_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput17 la_data_in[5] net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput28 la_oenb[15] net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_10_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput39 la_oenb[9] net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_42_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1437__A2 _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1984_ _1199_ _0414_ _0416_ _0055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2605_ u1.row_limit\[3\] _0877_ u1.row_limit\[2\] _0881_ _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__3100__CLK clknet_leaf_29_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2536_ _0380_ _0832_ _0833_ spi_data_crossing\[10\].data_sync _0836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3250__CLK clknet_leaf_8_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2467_ u1.ordering_timer\[26\] _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1418_ _1040_ u0.cmd\[30\] _1042_ _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_29_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2173__I0 _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2398_ _1096_ u1.ordering_timer\[14\] _0693_ _0722_ _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__2468__A4 _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2625__A1 net217 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1428__A2 u1.ordering_complete\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3019_ _0161_ clknet_leaf_13_clock u1.ordering_timer\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_25_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2968__CLK clknet_leaf_22_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2616__A1 _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1419__A2 control_trigger vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2092__A2 _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2219__I1 u1.row_col_select\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3123__CLK clknet_leaf_36_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2124__I u1.ordering_complete\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2060__S _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2321_ _0626_ _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2252_ _1095_ _0588_ _0590_ _0593_ _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2183_ _0461_ u1.inverter_select\[2\] _0540_ _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_38_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1658__A2 _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2743__B u1.timer\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2386__A3 _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1967_ _0396_ _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1898_ _0353_ _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2519_ _0825_ _0181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2689__A4 _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input31_I la_oenb[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1821__A2 u0.cmd\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2145__S _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3187__D _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold6 u0.mem_write_n\[5\] net248 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_43_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1958__I _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2870_ _0027_ clknet_leaf_14_clock u1.col_sel\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1821_ u0.cmd\[28\] u0.cmd\[29\] _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3097__D _0231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1752_ _1367_ u1.ccr0\[3\] _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1683_ u1.timer\[13\] _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3019__CLK clknet_leaf_13_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3284_ net100 net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2304_ _0613_ _0639_ _0640_ _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2235_ _1120_ _0570_ _0573_ _0576_ _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__2828__A1 net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3169__CLK clknet_leaf_7_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2166_ _0318_ _0530_ _0533_ _0120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_38_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2097_ _0488_ _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_22_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2999_ _0141_ clknet_leaf_18_clock u1.row_col_select\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2367__I0 u1.ordering_complete\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_21_clock_I clknet_2_3__leaf_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2648__B _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2819__A1 _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2295__A2 _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2020_ u1.ccr1\[21\] _0368_ _0432_ _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_36_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2922_ _0064_ clknet_leaf_2_clock u1.ccr1\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1797__A1 _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2853_ u0.cmd\[9\] clknet_leaf_16_clock net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2784_ _0393_ _0394_ _0351_ _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_1804_ u1.timer\[22\] _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1735_ u1.ccr0\[31\] _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1666_ _1190_ _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1597_ u1.ccr1\[2\] _1215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1721__A1 _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3267_ net86 net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2218_ _0562_ _0143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3198_ _0268_ clknet_leaf_23_clock u1.ccr0\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2149_ u1.row_limit\[4\] _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_26_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1788__A1 _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2650__C _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1520_ _1144_ _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1451_ u1.ordering_timer\[29\] _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_49_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3121_ spi_data_crossing\[1\].A clknet_leaf_35_clock spi_data_crossing\[1\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2851__CLK clknet_leaf_15_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3052_ _0194_ clknet_leaf_5_clock u0.cmd\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2259__A2 _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2003_ _0347_ _0395_ _0351_ _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_24_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2307__I _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3207__CLK clknet_leaf_35_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2431__A2 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2905_ _0047_ clknet_leaf_0_clock u1.ccr0\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2836_ net271 clknet_leaf_10_clock net208 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2767_ net11 _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2698_ _1248_ _0954_ _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1718_ _1233_ u1.ccr0\[21\] u1.ccr0\[20\] _1224_ _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1649_ u1.timer\[8\] _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_8_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2498__A2 _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1458__B1 _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output100_I net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2422__A2 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2874__CLK clknet_leaf_16_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2489__A2 _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2661__A2 _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2127__I u1.ordering_complete\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2413__A2 _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1966__I u0.cmd\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2063__S _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout229_I net233 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2621_ _0890_ _0895_ _0896_ _0212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__2177__A1 net218 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput105 net105 data_out_left[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput116 net116 data_out_right[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_2552_ _0819_ _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput127 net127 inverter_select[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_1503_ u1.ordering_timer\[3\] _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_5_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput149 net149 io_driver_io_oeb[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput138 net138 io_driver_io_oeb[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_12_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2483_ _0796_ _0791_ _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1434_ u1.ordering_timer\[16\] _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_28_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3104_ _0238_ clknet_leaf_30_clock u1.timer\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3035_ _0177_ clknet_leaf_22_clock u1.ordering_timer\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2101__A1 _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2652__A2 _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1860__C2 _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2819_ _1310_ _1025_ _1033_ _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input61_I spi_data[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2897__CLK clknet_leaf_2_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2340__A1 u1.ordering_complete\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2656__B _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2643__A2 _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput18 la_data_in[6] net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_7_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput29 la_oenb[16] net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__2159__A1 _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3052__CLK clknet_leaf_5_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2398__A1 _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1983_ _0373_ _0412_ _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2604_ u1.row_limit\[2\] _0881_ u1.row_limit\[1\] _0878_ _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2535_ _0835_ _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2466_ _0782_ _0171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1417_ _1041_ _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2173__I1 u1.col_limit\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2397_ _1068_ _1059_ _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_29_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3018_ _0160_ clknet_leaf_13_clock u1.ordering_timer\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_25_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2389__A1 u1.ordering_complete\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3075__CLK clknet_leaf_11_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2912__CLK clknet_leaf_24_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_16_clock_I clknet_2_3__leaf_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1465__B _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2140__I _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2320_ u1.ordering_timer\[8\] _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2251_ _1083_ _0592_ _1074_ _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2304__A1 _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2182_ _0542_ _0127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_19_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1966_ u0.cmd\[2\] _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3098__CLK clknet_leaf_27_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1897_ _0352_ _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2050__I _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2518_ _0364_ _0818_ _0821_ spi_data_crossing\[3\].data_sync _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2449_ _0767_ _0169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2935__CLK clknet_leaf_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input24_I la_oenb[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2782__A1 _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2534__B2 spi_data_crossing\[9\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2534__A1 _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold7 u1.output_active net249 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_48_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3240__CLK clknet_leaf_7_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1820_ _1040_ _0295_ u0.update_cmd _0022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_30_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2071__S _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1751_ _1367_ u1.ccr0\[3\] u1.ccr0\[2\] _1204_ _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1682_ _1293_ u1.ccr0\[9\] _1294_ _1298_ _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_48_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2958__CLK clknet_leaf_20_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2303_ u1.ordering_complete\[5\] _0630_ _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3283_ net99 net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2234_ _1114_ _0575_ _1108_ _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2165_ _0356_ _0531_ _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_22_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2096_ _0487_ _0454_ _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2998_ _0140_ clknet_leaf_18_clock u1.row_col_select\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1567__A2 _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1949_ net219 _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2764__A1 _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1811__I0 net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2516__B2 spi_data_crossing\[2\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2516__A1 _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3113__CLK clknet_leaf_34_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1552__C _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output130_I net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1730__A2 u1.ccr0\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2066__S _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2921_ _0063_ clknet_leaf_29_clock u1.ccr1\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1797__A2 u1.timer\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2852_ u0.cmd\[8\] clknet_leaf_16_clock net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1803_ _1327_ _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2783_ u1.ccr0\[0\] _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1734_ u1.timer\[31\] _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2761__A4 _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1665_ u1.ccr0\[5\] _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1596_ u1.timer\[3\] _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3266_ net85 net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1721__A2 u1.ccr0\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2217_ _0474_ u1.row_col_select\[7\] _0558_ _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3197_ _0267_ clknet_leaf_23_clock u1.ccr0\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2148_ _0520_ _0115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2079_ u0.cmd\[9\] _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1788__A2 _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2752__A4 _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3009__CLK clknet_leaf_16_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3159__CLK clknet_leaf_6_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1951__A2 _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1450_ _1071_ u1.ordering_complete\[28\] _1072_ u1.ordering_complete\[27\] _1074_
+ _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_45_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3120_ net51 net229 spi_data_crossing\[1\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3051_ _0193_ clknet_leaf_1_clock u0.cmd\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2002_ _1252_ _0405_ _0426_ _0063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2904_ _0046_ clknet_leaf_36_clock u1.ccr0\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2835_ u1.row_sel\[3\] clknet_leaf_10_clock net207 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2719__A1 _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2766_ _1001_ net30 _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2697_ _0951_ _0955_ _0956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1717_ _1236_ u1.ccr0\[17\] u1.ccr0\[16\] _1237_ _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__1942__A2 _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1648_ _1260_ _1265_ _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_28_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1579_ u1.ccr1\[4\] _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3249_ net248 clknet_leaf_10_clock net187 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1458__B2 _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2430__I0 u1.ordering_complete\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1697__A1 _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2620_ u1.row_sel\[1\] _0892_ u1.row_sel\[2\] _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput106 net106 data_out_left[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_2551_ _0844_ _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xoutput117 net117 data_out_right[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_47_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput128 net128 inverter_select[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_1502_ _1123_ _1126_ _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2482_ _1071_ _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput139 net139 io_driver_io_oeb[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_1433_ u1.ordering_complete\[19\] _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_3_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3103_ _0237_ clknet_leaf_32_clock u1.timer\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3034_ _0176_ clknet_leaf_22_clock u1.ordering_timer\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2101__A2 _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2818_ u0.cmd\[12\] _1029_ _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2168__A2 _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1892__I u0.cmd\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2749_ _1410_ _0990_ _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input54_I spi_data[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2002__B _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2340__A2 _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2391__C _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1603__A1 _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput19 la_data_in[7] net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_11_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2841__CLK clknet_leaf_15_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2159__A2 _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2991__CLK clknet_leaf_17_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_12_clock_I clknet_2_1__leaf_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1977__I _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2074__S _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout241_I net242 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2398__A2 u1.ordering_timer\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1982_ _1200_ _0414_ _0415_ _0054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2603_ u1.row_sel\[2\] _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2601__I u1.row_sel\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2534_ _0377_ _0832_ _0833_ spi_data_crossing\[9\].data_sync _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2465_ _0773_ _0754_ _0761_ _0781_ _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2396_ _0708_ _0712_ _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1416_ reset_n_sync\[1\] reset_n_sync\[0\] reset_n _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__2322__A2 _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2086__A1 _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2048__I _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3017_ _0159_ clknet_leaf_13_clock u1.ordering_timer\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_25_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2389__A2 _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2864__CLK clknet_leaf_4_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2511__I _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output160_I net160 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2001__A1 _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2250_ _1077_ _0591_ _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2181_ _0357_ u1.inverter_select\[1\] _0540_ _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_38_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1512__B1 _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2887__CLK clknet_leaf_8_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1815__A1 net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1500__I u1.ordering_timer\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1965_ _0402_ _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2240__A1 _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1896_ _0347_ _0348_ _0351_ _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2517_ _0824_ _0180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2448_ _0760_ _0754_ _0761_ _0766_ _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_9_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2379_ u1.ordering_complete\[15\] _0705_ _0609_ _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_29_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input17_I la_data_in[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3042__CLK clknet_leaf_3_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2241__I u1.ordering_timer\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output85_I net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3192__CLK clknet_leaf_30_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold8 control_trigger net250 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_16_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2470__A1 _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1750_ _1214_ _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_8_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1681_ _1295_ _1296_ _1297_ _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_7_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2302_ _0636_ _0638_ _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1733__B1 u1.ccr0\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3282_ net98 net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input9_I la_data_in[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2233_ _1117_ _0574_ _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2164_ _0321_ _0530_ _0532_ _0119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_26_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2095_ _0347_ _0394_ _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_19_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3065__CLK clknet_leaf_6_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2461__A1 _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2997_ _0139_ clknet_leaf_16_clock u1.row_col_select\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1948_ _1353_ _0362_ _0389_ _0046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1879_ u1.col_sel\[3\] _0336_ _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1811__I1 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2902__CLK clknet_leaf_36_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2452__A1 u1.ordering_complete\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2755__A2 _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3088__CLK clknet_leaf_29_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2920_ _0062_ clknet_leaf_28_clock u1.ccr1\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2851_ u0.cmd\[7\] clknet_leaf_15_clock net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2782_ _1009_ net39 _0260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1802_ _0281_ _1322_ _0282_ _0283_ _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__2925__CLK clknet_leaf_30_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2746__A2 _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1733_ _1173_ u1.ccr0\[28\] u1.ccr0\[27\] _1349_ _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_15_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2810__S _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1664_ u1.ccr0\[6\] _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1706__B1 _1320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1595_ u1.ccr1\[3\] _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3265_ net84 net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2216_ _0561_ _0142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3196_ _0266_ clknet_leaf_24_clock u1.ccr0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2147_ _0464_ u1.row_limit\[3\] _0515_ _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2682__A1 _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2078_ _0477_ _0088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2056__I _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3230__CLK clknet_leaf_17_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2948__CLK clknet_leaf_12_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2425__A1 u1.ordering_timer\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2841__D u1.col_sel\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1754__B _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3050_ _0192_ clknet_leaf_1_clock u0.cmd\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2001_ _0390_ _0398_ _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3260__I clknet_leaf_10_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2077__S _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2664__A1 _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2416__A1 _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2903_ _0045_ clknet_leaf_36_clock u1.ccr0\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2834_ u1.row_sel\[2\] clknet_leaf_9_clock net206 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3103__CLK clknet_leaf_32_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2765_ net12 _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2696_ _1293_ _1267_ _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1716_ _1330_ _1332_ _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3253__CLK clknet_leaf_9_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1647_ _1261_ _1262_ _1264_ _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1578_ u1.ccr1\[5\] _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_41_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3248_ net247 clknet_leaf_9_clock net186 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3179_ spi_data_crossing\[30\].A clknet_leaf_6_clock spi_data_crossing\[30\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1458__A2 _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2655__A1 u1.ccr1\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2407__A1 _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2194__I0 _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1697__A2 u1.ccr0\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2646__A1 _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1449__A2 _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput107 net107 data_out_left[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_2550_ _0816_ _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xoutput118 net118 data_out_right[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__3255__I clknet_leaf_9_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput129 net129 inverter_select[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_1501_ _1124_ u1.ordering_complete\[7\] _1125_ u1.ordering_complete\[6\] _1126_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2481_ _1093_ _0710_ _0795_ _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1432_ _1052_ _1053_ _1056_ _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__2185__I0 _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3102_ _0236_ clknet_leaf_28_clock u1.timer\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2637__A1 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3033_ _0175_ clknet_leaf_22_clock u1.ordering_timer\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1860__A2 u1.col_limit\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2762__C _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2817_ _1031_ _1025_ _1032_ _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2748_ _0983_ _0989_ _0990_ _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2679_ _1287_ _0941_ _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_28_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input47_I spi_data[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3149__CLK clknet_leaf_1_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output203_I net203 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2619__A1 u1.row_sel\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1981_ _0370_ _0412_ _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2602_ u1.row_limit\[1\] _0878_ u1.row_limit\[0\] _0879_ _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2533_ _0834_ _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_29_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2464_ u1.ordering_complete\[25\] _0779_ _0780_ _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_9_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1415_ u0.cmd\[31\] _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2395_ _0612_ _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_25_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1530__A1 _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2086__A2 _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3016_ _0158_ clknet_leaf_14_clock u1.ordering_timer\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_25_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3100__D _0234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1824__A2 _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2180_ _0541_ _0126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1512__A1 _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1964_ _0397_ _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2240__A2 _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1895_ _0349_ _0350_ _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2379__I0 u1.ordering_complete\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2516_ _0361_ _0818_ _0821_ spi_data_crossing\[2\].data_sync _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2447_ _1054_ _0720_ _0765_ _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1751__B2 _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2059__I _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2378_ _0703_ _0704_ _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_25_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1898__I _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1806__A2 _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2981__CLK clknet_leaf_16_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2231__A2 u1.ordering_complete\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold9 u0.mem_write_n\[1\] net251 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_43_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2844__D u0.cmd\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1680_ _1269_ u1.ccr0\[11\] _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1981__A1 _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2301_ _1121_ _0637_ _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1733__A1 _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3263__I clknet_leaf_10_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3281_ net97 net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2854__CLK clknet_leaf_16_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2232_ _1109_ _1110_ _1111_ u1.ordering_complete\[8\] _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2163_ _0345_ _0531_ _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2808__S _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2094_ _1097_ _0458_ _0486_ _0095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1511__I u1.ordering_timer\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2996_ _0138_ clknet_leaf_16_clock u1.row_col_select\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1947_ _0388_ _0384_ _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1878_ u1.col_sel\[3\] _0336_ _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_31_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2517__I _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1421__I u1.ordering_timer\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2452__A2 _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2877__CLK clknet_leaf_12_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2850_ u0.cmd\[6\] clknet_leaf_15_clock net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1801_ u1.timer\[16\] _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3258__I clknet_leaf_9_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2162__I _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2781_ net21 _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_12_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1732_ _1177_ _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_7_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1663_ _1188_ _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1594_ u0.timer_enable _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1706__A1 _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1706__B2 _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3264_ net83 net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2215_ _0471_ u1.row_col_select\[6\] _0558_ _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3032__CLK clknet_leaf_21_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3195_ _0265_ clknet_leaf_23_clock u1.ccr0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2146_ _0519_ _0114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2077_ _0476_ _1112_ _0472_ _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2337__I _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3182__CLK clknet_leaf_32_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2979_ _0121_ clknet_leaf_14_clock u1.col_limit\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2183__S _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1936__A1 _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3055__CLK clknet_leaf_5_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2000_ _1253_ _0421_ _0425_ _0062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_49_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2902_ _0044_ clknet_leaf_36_clock u1.ccr0\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2833_ net293 clknet_leaf_10_clock net205 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2764_ _1351_ _0999_ _1000_ _0934_ _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__2719__A3 _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1715_ _1229_ u1.ccr0\[22\] _1331_ _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2695_ _0946_ _0953_ _0954_ _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_6_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1646_ _1263_ u1.timer\[13\] _1261_ u1.timer\[12\] _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_28_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1577_ u1.ccr1\[7\] _1193_ u1.ccr1\[4\] _1194_ _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_28_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3247_ net255 clknet_leaf_8_clock net185 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2104__A1 _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2495__C _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3178_ net63 net237 spi_data_crossing\[30\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2129_ u0.cmd\[11\] _0509_ _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3078__CLK clknet_leaf_9_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2530__I _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2915__CLK clknet_leaf_26_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2646__A2 _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2852__D u0.cmd\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1909__A1 _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput119 net119 data_out_right[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput108 net108 data_out_left[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_1500_ u1.ordering_timer\[6\] _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2480_ _0793_ _0794_ _0604_ _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1431_ _1050_ u1.ordering_complete\[20\] _1055_ _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2334__A1 _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput90 net90 col_select_right[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_3101_ _0235_ clknet_leaf_28_clock u1.timer\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3271__I net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3032_ _0174_ clknet_leaf_21_clock u1.ordering_timer\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2270__B1 _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3220__CLK clknet_leaf_17_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2816_ net223 _1029_ _1032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2747_ _1411_ _0988_ _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2678_ _1287_ _0941_ _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1629_ u1.ccr1\[9\] _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2325__A1 _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2938__CLK clknet_leaf_12_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2800__A2 _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2564__A1 u0.cmd\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2260__I _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2316__A1 u1.ordering_complete\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2847__D net288 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2619__A2 u1.row_sel\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3243__CLK clknet_leaf_7_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1980_ _0402_ _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_fanout227_I net229 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3266__I net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2601_ u1.row_sel\[0\] _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_9_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2532_ _0375_ _0832_ _0833_ spi_data_crossing\[8\].data_sync _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2463_ _0607_ _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_29_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2394_ _0626_ _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3015_ _0157_ clknet_leaf_14_clock u1.ordering_timer\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2345__I _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2546__B2 spi_data_crossing\[14\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2546__A1 _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3116__CLK clknet_leaf_36_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1424__I u1.ordering_timer\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output146_I net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2255__I _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_hold48_I u0.cmd\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1512__A2 u1.ordering_complete\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2473__B1 _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1963_ _0401_ _0049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1894_ u0.write_config_n u0.cmd\[18\] u0.cmd\[21\] u0.cmd\[20\] _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__2776__A1 _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2240__A3 _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1509__I u1.ordering_complete\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2528__B2 spi_data_crossing\[7\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2528__A1 _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3139__CLK clknet_leaf_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2515_ _0823_ _0179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2446_ _0756_ _0763_ _0764_ _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__1751__A2 u1.ccr0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_2_0__f_clock clknet_0_clock clknet_2_0__leaf_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_2377_ _0698_ _0694_ _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2860__D net249 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1430__A1 u1.ordering_timer\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3280_ net96 net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2300_ _0625_ _0628_ _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1733__A2 u1.ccr0\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2231_ _0571_ u1.ordering_complete\[15\] _1099_ _0572_ _0573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2162_ _0528_ _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2093_ net219 _0480_ _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_4_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2995_ _0137_ clknet_leaf_16_clock u1.row_col_select\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1946_ net220 _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1877_ _0330_ _0336_ _0337_ _0027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_31_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1972__A2 _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2221__I0 _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2429_ _1049_ _0745_ _0749_ _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1903__S _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input22_I la_oenb[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output109_I net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1715__A2 u1.ccr0\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_2_3__f_clock_I clknet_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2855__D net223 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1612__I u1.timer\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1800_ u1.timer\[17\] _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2780_ _1008_ net23 _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_12_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1731_ _1180_ u1.ccr0\[26\] u1.ccr0\[25\] _1164_ _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_15_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1662_ _1279_ u1.ccr1_flag vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3274__I net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1706__A2 _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1593_ _1205_ _1210_ _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3263_ clknet_leaf_10_clock net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2214_ _0560_ _0141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2971__CLK clknet_leaf_11_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3194_ _0264_ clknet_leaf_30_clock u1.ccr0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2145_ _0461_ u1.row_limit\[2\] _0515_ _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_27_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2076_ u0.cmd\[8\] _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2978_ _0120_ clknet_leaf_11_clock u1.col_limit\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1929_ _0376_ _0040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1945__A2 _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2464__S _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2263__I _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1633__B2 _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2844__CLK clknet_leaf_15_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1936__A2 _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2994__CLK clknet_leaf_16_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1607__I u1.ccr1\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2664__A3 _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1872__A1 _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2901_ _0043_ clknet_leaf_34_clock u1.ccr0\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1624__A1 u1.ccr1\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3269__I net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2832_ net292 clknet_leaf_10_clock net204 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2763_ _1351_ _0999_ _1000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1714_ _1327_ _1328_ _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2694_ _1250_ _0951_ _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1645_ u1.ccr1\[13\] _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1576_ u1.timer\[4\] _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_8_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3246_ net256 clknet_leaf_8_clock net184 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2104__A2 _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3177_ spi_data_crossing\[29\].A clknet_leaf_7_clock spi_data_crossing\[29\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2128_ _0491_ _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2059_ _0407_ _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2867__CLK clknet_leaf_32_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2031__A1 _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1909__A2 _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3022__CLK clknet_leaf_30_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput109 net109 data_out_left[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_5_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3172__CLK net240 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1430_ u1.ordering_timer\[23\] _1054_ _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2334__A2 _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput91 net91 col_select_right[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput80 net80 clock_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
XANTENNA__1542__B1 _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3100_ _0234_ clknet_leaf_29_clock u1.timer\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3031_ _0173_ clknet_leaf_24_clock u1.ordering_timer\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2815_ u1.ccr0\[11\] _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2746_ _1411_ _0988_ _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2022__A1 _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2677_ _0937_ _0940_ _0941_ _0223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1628_ _1235_ _1245_ _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2325__A2 _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1559_ u1.timer\[27\] _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3229_ net280 clknet_leaf_18_clock net199 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1836__A1 _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3045__CLK clknet_leaf_1_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2541__I _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3195__CLK clknet_leaf_23_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2316__A2 _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2863__D net250 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2252__A1 _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2600_ u1.row_sel\[1\] _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2531_ _0820_ _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2462_ _0773_ _0778_ _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__3282__I net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2393_ _0708_ _0710_ _0718_ _0162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3014_ _0156_ clknet_leaf_21_clock u1.ordering_timer\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3068__CLK clknet_leaf_4_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2491__A1 _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2491__B2 _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2905__CLK clknet_leaf_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2729_ _0281_ _1322_ _0974_ _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA_input52_I spi_data[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1506__B1 _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1705__I _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1440__I u1.ordering_timer\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2234__A1 _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2858__D net220 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1899__I1 _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3210__CLK clknet_leaf_35_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2225__A1 _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2928__CLK clknet_leaf_31_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1962_ u1.ccr1\[1\] _0400_ _0398_ _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3277__I net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1893_ net218 _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_18_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2514_ _0400_ _0818_ _0821_ spi_data_crossing\[1\].data_sync _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2445_ _0760_ _0753_ _0749_ _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__2130__B _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2376_ _1096_ _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3233__CLK clknet_leaf_17_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1435__I u1.ordering_complete\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2266__I _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1718__B1 u1.ccr0\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2230_ _1102_ _1106_ _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2161_ _0529_ _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2694__A1 _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2092_ _1098_ _0458_ _0485_ _0094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2446__A1 _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3212__D _0002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2994_ _0136_ clknet_leaf_16_clock u1.row_col_select\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2461__A4 _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1945_ _1357_ _0379_ _0387_ _0045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3106__CLK clknet_leaf_31_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1876_ _0317_ _0333_ net225 _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_27_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2428_ _0748_ _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2359_ _0670_ _0686_ _0688_ _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2437__A1 u1.ordering_complete\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input15_I la_data_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3122__D net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1660__A2 _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3129__CLK clknet_leaf_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1730_ _1164_ u1.ccr0\[25\] u1.ccr0\[24\] _1166_ _1346_ _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_1661_ _1187_ _1222_ _1278_ _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__1784__B _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1592_ _1207_ u1.ccr1\[0\] u1.ccr1\[1\] _1209_ _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1962__I0 u1.ccr1\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3262_ clknet_leaf_10_clock net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2213_ _0368_ u1.row_col_select\[5\] _0558_ _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_26_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input7_I la_data_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3193_ _0263_ clknet_leaf_30_clock u1.ccr0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2144_ _0518_ _0113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2075_ _0475_ _0087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2419__A1 _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2977_ _0119_ clknet_leaf_11_clock u1.col_limit\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1928_ u1.ccr0\[24\] _0375_ _0359_ _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1859_ net226 _0321_ u1.col_sel\[1\] _0318_ _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2830__A1 net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1633__A2 _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2649__A1 _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1872__A2 _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2900_ _0042_ clknet_leaf_34_clock u1.ccr0\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1624__A2 _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2831_ _1039_ _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2762_ _1167_ _0998_ _0999_ _0934_ _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__3285__I net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1713_ _1327_ _1328_ _1329_ u1.timer\[22\] _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2693_ _1250_ _0951_ _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2188__I0 _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1644_ u1.timer\[12\] _1262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1575_ u1.timer\[7\] _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3245_ net251 clknet_leaf_8_clock net183 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3176_ net61 net238 spi_data_crossing\[29\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2127_ u1.ordering_complete\[27\] _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2058_ _0463_ _0082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2576__B1 _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2179__I0 _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output169_I net169 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2803__A1 _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2961__CLK clknet_leaf_21_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2031__A2 _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput92 net92 col_select_right[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput81 net81 clock_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
XANTENNA__1542__B2 _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2449__I _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3030_ _0172_ clknet_leaf_24_clock u1.ordering_timer\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3220__D net281 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2270__A2 _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2814_ _1296_ _1025_ _1030_ _0271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2745_ _0983_ _0987_ _0988_ _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__2022__A2 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2676_ u1.timer\[0\] u1.timer\[1\] u1.timer\[3\] u1.timer\[2\] _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__1781__A1 _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1627_ _1238_ _1244_ _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_28_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1533__A1 _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1558_ u1.ccr1\[27\] _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1489_ u1.ordering_timer\[11\] _1104_ u1.ordering_timer\[10\] _1113_ _1114_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2834__CLK clknet_leaf_9_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3228_ net263 clknet_leaf_17_clock net198 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1836__A2 _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3159_ spi_data_crossing\[20\].A clknet_leaf_6_clock spi_data_crossing\[20\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2984__CLK clknet_leaf_18_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1524__A1 u0.cmd\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2721__B1 _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1901__I u0.cmd\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2530_ _0817_ _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2461_ _1085_ _0760_ _0753_ _0777_ _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_5_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2857__CLK clknet_leaf_15_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2400__C _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2392_ _0329_ _0717_ _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3013_ _0155_ clknet_leaf_19_clock u1.ordering_timer\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2728_ _0281_ _0976_ _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2659_ _1187_ _0926_ _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1506__B2 u1.ordering_complete\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input45_I spi_data[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3012__CLK clknet_leaf_19_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output201_I net201 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3162__CLK net239 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1993__A1 _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1631__I u1.ccr1\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2473__A2 _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2225__A2 _1140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1961_ u0.cmd\[1\] _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1892_ u0.cmd\[17\] _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout232_I net233 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1984__A1 _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2513_ _0822_ _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2444_ _1046_ _0762_ _0763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2375_ _0702_ _0160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3035__CLK clknet_leaf_22_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3185__CLK clknet_leaf_33_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1718__B2 _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1718__A1 _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3058__CLK clknet_leaf_6_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2391__A1 _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2160_ _0528_ _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_26_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2091_ net220 _0480_ _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_47_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2993_ _0135_ clknet_leaf_18_clock u1.inverter_select\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1944_ _0386_ _0384_ _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1875_ _0317_ net225 _0333_ _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2427_ _0583_ u1.ordering_timer\[18\] _0723_ _0747_ _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_9_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2358_ u1.ordering_complete\[12\] _0687_ _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_42_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2289_ _0626_ _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2437__A2 _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3200__CLK clknet_leaf_31_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1446__I u1.ordering_timer\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2373__A1 _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2918__CLK clknet_leaf_27_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2125__A1 u0.cmd\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2676__A2 u1.timer\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1939__A1 _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1660_ _1246_ _1277_ _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1591_ _1208_ _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_4_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1962__I1 _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3261_ clknet_leaf_10_clock net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2212_ _0559_ _0140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3192_ _0262_ clknet_leaf_30_clock u1.ccr0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2187__I _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2143_ _0357_ u1.row_limit\[1\] _0516_ _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2074_ _0474_ u1.ordering_complete\[7\] _0472_ _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2419__A2 _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3223__CLK clknet_leaf_17_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2976_ _0118_ clknet_leaf_11_clock u1.row_limit\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1975__B _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1927_ u0.cmd\[8\] _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1858_ u1.col_limit\[0\] _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_11_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1789_ _1289_ _1280_ _1283_ _1287_ _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_44_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2658__A2 _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2097__I _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3133__D spi_data_crossing\[7\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2594__A1 _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2346__A1 _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold16_I u0.cmd\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2890__CLK clknet_leaf_3_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3246__CLK clknet_leaf_8_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2735__I _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2830_ net14 net32 _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_32_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2761_ u1.timer\[30\] _0996_ _1413_ _0993_ _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_1712_ u1.ccr0\[22\] _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2692_ _0946_ _0951_ _0952_ _0227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1643_ u1.ccr1\[12\] _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_clkbuf_0_clock_I clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1574_ u1.ccr1\[6\] _1189_ u1.ccr1\[5\] _1191_ _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3244_ net252 clknet_leaf_8_clock net182 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3175_ spi_data_crossing\[28\].A clknet_leaf_7_clock spi_data_crossing\[28\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2126_ _0506_ _0502_ _0507_ _0106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_39_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2057_ _0461_ u1.ordering_complete\[2\] _0462_ _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2959_ _0101_ clknet_leaf_20_clock u1.ordering_complete\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3119__CLK clknet_leaf_35_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_6_clock_I clknet_2_1__leaf_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2500__A1 u1.ordering_timer\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2803__A2 _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput82 net82 clock_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
Xoutput93 net93 col_select_right[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_1_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3296__I net162 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2813_ net224 _1029_ _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2558__A1 u0.cmd\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2744_ u1.timer\[24\] _1327_ _0286_ _0981_ _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2675_ _1214_ _0938_ _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1626_ _1241_ _1242_ _1243_ _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1557_ _1172_ _1174_ _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__1533__A2 u0.cmd\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2730__A1 _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1488_ u1.ordering_complete\[10\] _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3227_ net274 clknet_leaf_17_clock net197 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3158_ net52 net235 spi_data_crossing\[20\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2375__I _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2109_ _1058_ _0490_ _0497_ _0099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_39_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3089_ _0223_ clknet_leaf_29_clock u1.timer\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2246__B1 _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output181_I net181 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1454__I u1.ordering_complete\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2721__A1 _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3091__CLK clknet_leaf_25_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2234__B _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2460_ _1064_ _0728_ _0776_ _0746_ _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__1763__A2 _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1515__A2 _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2391_ _0711_ _0713_ _0715_ _0716_ _0717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__2712__A1 _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3012_ _0154_ clknet_leaf_19_clock u1.ordering_timer\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1539__I _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2727_ _0968_ _0975_ _0976_ _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__1754__A2 u1.ccr0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2658_ _1246_ _0918_ _0925_ _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1506__A2 u1.ordering_complete\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2589_ _0868_ _0208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2703__A1 _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1609_ _1225_ u1.timer\[23\] _1226_ u1.timer\[22\] _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_47_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input38_I la_oenb[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2951__CLK clknet_leaf_4_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1690__A1 _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1690__B2 _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1993__A2 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1960_ _0399_ _0048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1891_ u0.cmd\[16\] _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_35_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2512_ _0392_ _0818_ _0821_ spi_data_crossing\[0\].data_sync _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2974__CLK clknet_leaf_11_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2443_ _0753_ _0749_ _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2374_ _0698_ _0682_ _0691_ _0701_ _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_25_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_33_clock_I clknet_2_0__leaf_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1975__A2 _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2563__I _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2847__CLK clknet_leaf_10_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2215__I0 _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2997__CLK clknet_leaf_16_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1907__I u0.cmd\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold46_I u0.cmd\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2090_ _0484_ _0093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2446__A3 _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2992_ _0134_ clknet_leaf_18_clock u1.inverter_select\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1943_ net221 _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2206__I0 _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1874_ _0331_ _0335_ _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_31_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3002__CLK clknet_leaf_18_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2426_ _0746_ _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2134__A2 _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2357_ _0596_ _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2288_ _0600_ _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2383__I _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1928__S _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1948__A2 _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1727__I u1.ccr0\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2125__A2 _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1462__I u1.ordering_timer\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3025__CLK clknet_leaf_20_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1939__A2 _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3175__CLK clknet_leaf_7_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1590_ u1.timer\[1\] _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2364__A2 _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3260_ clknet_leaf_10_clock net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2211_ _0366_ u1.row_col_select\[4\] _0558_ _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3191_ _0261_ clknet_leaf_23_clock u1.ccr0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1875__A1 _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2142_ _0517_ _0112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2073_ u0.cmd\[7\] _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3299__I net165 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2975_ _0117_ clknet_leaf_11_clock u1.row_limit\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2052__A1 _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1926_ _1328_ _0360_ _0374_ _0039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1857_ _0317_ _0318_ net225 _0319_ _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1547__I u1.timer\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2355__A2 _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1788_ _1256_ _1257_ _1258_ _1404_ _1405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__2107__A2 _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2409_ _0728_ _0710_ _0732_ _0164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input20_I la_data_in[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output107_I net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2291__A1 _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3048__CLK clknet_leaf_5_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_2_clock_I clknet_2_0__leaf_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3198__CLK clknet_leaf_23_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1457__I u1.ordering_timer\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2346__A2 _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2288__I _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1857__A1 _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1920__I u0.cmd\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2760_ _0996_ _0995_ _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1711_ u1.ccr0\[23\] _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2691_ _1289_ _0948_ _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_32_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1642_ _1255_ _1259_ _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1573_ _1190_ _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3312_ net209 net215 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3243_ net286 clknet_leaf_7_clock net171 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3234__D u0.cmd\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3174_ net60 net240 spi_data_crossing\[28\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2125_ u0.cmd\[10\] _0495_ _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2056_ _0455_ _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_2_2__f_clock_I clknet_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2958_ _0100_ clknet_leaf_20_clock u1.ordering_complete\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2908__CLK clknet_leaf_22_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2576__A2 _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1909_ _0361_ _0362_ _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2889_ net279 clknet_leaf_3_clock u1.u1.impulse_gen\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input68_I spi_data[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1839__A1 _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2016__A1 _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1790__A3 _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput83 net83 col_select_left[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput94 net94 col_select_right[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_27_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3213__CLK clknet_leaf_32_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2812_ _1011_ _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2743_ _0285_ _0985_ u1.timer\[24\] _0987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2674_ _0937_ _0938_ _0939_ _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__1825__I u0.cmd\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1625_ u1.ccr1\[16\] _1237_ _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1556_ u1.ccr1\[29\] _1168_ u1.ccr1\[28\] _1173_ _1174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__1533__A3 _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1487_ u1.ordering_complete\[8\] _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3226_ net283 clknet_leaf_16_clock net196 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_2_3__f_clock clknet_0_clock clknet_2_3__leaf_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3157_ spi_data_crossing\[19\].A clknet_leaf_5_clock spi_data_crossing\[19\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2494__A1 u1.ordering_timer\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2108_ _0407_ _0495_ _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_36_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3088_ _0222_ clknet_leaf_29_clock u1.timer\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2246__B2 _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2246__A1 _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2039_ _0449_ _0077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2880__CLK clknet_leaf_8_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_28_clock_I clknet_2_2__leaf_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3236__CLK clknet_leaf_7_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1735__I u1.ccr0\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2485__A1 u1.ordering_complete\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2237__A1 _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2007__S _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1748__B1 u1.ccr0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2888__D u1.ccr1_flag vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1645__I u1.ccr1\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2390_ _0601_ _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3011_ _0153_ clknet_leaf_19_clock u1.ordering_timer\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2476__A1 u1.ordering_timer\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2228__B2 _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3109__CLK clknet_leaf_31_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2400__A1 _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2726_ _1321_ _0282_ u1.timer\[16\] _0970_ _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_12_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2657_ _0919_ _1234_ _1235_ _0923_ _0924_ _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_1608_ u1.ccr1\[22\] _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2588_ u0.cmd\[30\] _0864_ _0865_ spi_data_crossing\[30\].data_sync _0868_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1539_ _1158_ _0011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3209_ _0001_ clknet_leaf_28_clock net161 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output99_I net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2630__A1 _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1890_ _0345_ _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout218_I u0.cmd\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2511_ _0820_ _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2442_ _0603_ _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2373_ _0670_ _0699_ _0700_ _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_29_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3081__CLK clknet_leaf_4_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2621__A1 _0890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2709_ _0958_ _0963_ _0964_ _0232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA_input50_I spi_data[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2688__A1 _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2612__A1 _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2020__S _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2991_ _0133_ clknet_leaf_17_clock u1.inverter_select\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1942_ _1358_ _0379_ _0385_ _0044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1873_ _0317_ _0333_ _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__2941__CLK clknet_leaf_14_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3237__D net218 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1833__I u0.cmd\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2425_ u1.ordering_timer\[21\] u1.ordering_timer\[20\] _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2356_ _0684_ _0685_ _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2287_ u1.ordering_timer\[4\] _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1884__A2 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2964__CLK clknet_leaf_24_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2364__A3 _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2210_ _0552_ _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_26_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3190_ _0260_ clknet_leaf_35_clock net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2141_ _0346_ u1.row_limit\[0\] _0516_ _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_26_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2072_ _0473_ _0086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2824__A1 net219 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2974_ _0116_ clknet_leaf_11_clock u1.row_limit\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1925_ _0373_ _0371_ _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2052__A2 _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1856_ u1.col_limit\[2\] _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1787_ _1311_ _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2837__CLK clknet_leaf_10_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2408_ _0329_ _0731_ _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2339_ u1.ordering_timer\[10\] _0665_ _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2115__I0 _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input13_I la_data_in[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2987__CLK clknet_leaf_18_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2291__A2 _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1473__I u1.ordering_complete\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold50 u1.row_sel\[0\] net292 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_21_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2806__A1 _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2034__A2 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1710_ u1.timer\[23\] _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2690_ _0950_ _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1641_ u1.ccr1\[15\] _1256_ u1.ccr1\[14\] _1257_ u1.ccr1\[13\] _1258_ _1259_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_6_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3311_ net208 net214 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1572_ u1.timer\[5\] _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3242_ net285 clknet_leaf_7_clock net170 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3173_ spi_data_crossing\[27\].A clknet_leaf_7_clock spi_data_crossing\[27\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input5_I la_data_in[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2124_ u1.ordering_complete\[26\] _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2055_ _0404_ _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1481__B1 _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2957_ _0099_ clknet_leaf_3_clock u1.ordering_complete\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2025__A2 _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2888_ u1.ccr1_flag clknet_leaf_3_clock u1.u1.impulse_gen\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1908_ _0353_ _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1839_ _0304_ _1153_ _0298_ _0020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_11_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1784__A1 _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3015__CLK clknet_leaf_14_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_24_clock_I clknet_2_2__leaf_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3165__CLK clknet_leaf_6_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2016__A2 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1790__A4 _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput84 net84 col_select_left[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput73 net73 clock_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
XFILLER_1_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput95 net95 data_out_left[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_1_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2811_ _1028_ _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2742_ _0285_ _0985_ _0986_ _0982_ _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_34_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2673_ _1206_ _1208_ _1203_ _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1624_ u1.ccr1\[17\] _1236_ _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1555_ u1.timer\[28\] _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3038__CLK clknet_leaf_3_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3225_ net273 clknet_leaf_17_clock net195 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1486_ u1.ordering_timer\[8\] _1111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3156_ net50 net235 spi_data_crossing\[19\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2494__A2 _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3188__CLK clknet_leaf_33_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2107_ _1067_ _0490_ _0496_ _0098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3087_ _0221_ clknet_leaf_29_clock u1.timer\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2038_ u1.ccr1\[29\] _0386_ _0443_ _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_35_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2246__A2 _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1757__A1 _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2113__S _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output167_I net167 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2485__A2 _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2582__I _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2237__A2 _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2796__I0 u1.ccr0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3010_ _0152_ clknet_leaf_19_clock u1.ordering_timer\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2725_ _1322_ _0974_ _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2656_ u1.ccr1\[23\] _1228_ _1227_ _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_12_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1607_ u1.ccr1\[23\] _1225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2587_ _0867_ _0207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1538_ u0.run_state\[3\] u0.run_state\[4\] _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__2667__I _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1571__I _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1469_ _1093_ u1.ordering_complete\[27\] _1087_ u1.ordering_complete\[26\] _1094_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_47_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3208_ _0278_ clknet_leaf_35_clock net158 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3139_ spi_data_crossing\[10\].A clknet_leaf_0_clock spi_data_crossing\[10\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1978__A1 _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3203__CLK clknet_leaf_23_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2458__A2 _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2018__S _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2510_ _0819_ _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2441_ u1.ordering_timer\[23\] _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2372_ u1.ordering_complete\[14\] _0687_ _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_29_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2870__CLK clknet_leaf_14_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3226__CLK clknet_leaf_16_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2621__A2 _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2708_ _1311_ _0961_ _0964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2639_ _0906_ _1270_ _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2137__A1 u0.cmd\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input43_I spi_data[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1476__I u1.ordering_timer\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2679__A2 _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2893__CLK clknet_leaf_2_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2100__I _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3249__CLK clknet_leaf_10_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2990_ _0132_ clknet_leaf_17_clock u1.inverter_select\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1941_ net222 _0384_ _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1872_ _0331_ _0333_ _0334_ _0025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_7_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2211__S _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2424_ u1.ordering_timer\[20\] _0736_ _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2355_ u1.ordering_timer\[12\] _0675_ _0677_ _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_28_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2010__I _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2286_ _0624_ _0149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_42_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2358__A1 u1.ordering_complete\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2597__A1 _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_19_clock_I clknet_2_3__leaf_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2349__A1 _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold51_I u1.row_sel\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1934__I net224 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3071__CLK clknet_leaf_9_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1875__A3 _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2140_ _0515_ _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2071_ _0471_ u1.ordering_complete\[6\] _0472_ _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2765__I net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2285__B1 _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2824__A2 _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2973_ _0115_ clknet_leaf_11_clock u1.row_limit\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2206__S _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2588__A1 u0.cmd\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1924_ u0.cmd\[7\] _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_33_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3248__D net247 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1855_ u1.col_limit\[1\] _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1786_ _1402_ _1144_ _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2060__I0 _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2407_ _0711_ _0729_ _0730_ _0716_ _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__2512__A1 _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2338_ _0612_ _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2512__B2 spi_data_crossing\[0\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2269_ u1.ordering_complete\[1\] _0606_ _0609_ _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2115__I1 u1.ordering_complete\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_20_clock_I clknet_2_3__leaf_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output197_I net197 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3094__CLK clknet_leaf_26_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1554__A2 _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2503__A1 _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold40 u1.inverter_select\[7\] net282 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_29_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold51 u1.row_sel\[1\] net293 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2931__CLK clknet_leaf_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2806__A2 _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1490__B2 _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2026__S _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3068__D _0023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1640_ u1.timer\[13\] _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1571_ _1188_ _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3310_ net207 net213 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2742__A1 _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3241_ net254 clknet_leaf_7_clock net169 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3172_ net59 net240 spi_data_crossing\[27\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2123_ _0505_ _0105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2054_ _1134_ _0457_ _0460_ _0081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_35_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1481__B2 u1.ordering_complete\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2956_ _0098_ clknet_leaf_3_clock u1.ordering_complete\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2887_ _0021_ clknet_leaf_8_clock u0.mem_write_n\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1907_ u0.cmd\[2\] _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1838_ _0299_ _1160_ _0302_ _0305_ _0019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_11_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1769_ _1375_ _1381_ _1383_ _1384_ _1385_ _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XTAP_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2954__CLK clknet_leaf_3_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1839__A3 _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1527__A2 _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1484__I u1.ordering_timer\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2724__A1 _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput85 net85 col_select_left[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput74 net74 clock_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
XFILLER_49_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput96 net96 data_out_left[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_27_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2810_ u1.ccr0\[9\] _0377_ _1013_ _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2741_ _0285_ _0985_ _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_8_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2672_ _1364_ _1363_ _1204_ _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__2977__CLK clknet_leaf_11_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1518__A2 _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1623_ _1239_ _1240_ _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1554_ u1.ccr1\[31\] _1171_ u1.ccr1\[30\] _1167_ _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1485_ u1.ordering_complete\[9\] _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3224_ net287 clknet_leaf_16_clock net194 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
.ends

